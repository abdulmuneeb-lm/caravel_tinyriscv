VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tinyriscv
  CLASS BLOCK ;
  FOREIGN tinyriscv ;
  ORIGIN 0.000 0.000 ;
  SIZE 1098.305 BY 1109.025 ;
  PIN int_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END int_i[0]
  PIN int_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 32.680 1098.305 33.280 ;
    END
  END int_i[1]
  PIN int_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END int_i[2]
  PIN int_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END int_i[3]
  PIN int_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.610 1105.025 281.890 1109.025 ;
    END
  END int_i[4]
  PIN int_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 1105.025 44.530 1109.025 ;
    END
  END int_i[5]
  PIN int_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 672.610 1105.025 672.890 1109.025 ;
    END
  END int_i[6]
  PIN int_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END int_i[7]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 934.810 1105.025 935.090 1109.025 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1015.770 0.000 1016.050 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 924.840 1098.305 925.440 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 857.530 0.000 857.810 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.370 1105.025 123.650 1109.025 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.490 1105.025 202.770 1109.025 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 405.320 1098.305 405.920 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.810 1105.025 544.090 1109.025 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 773.810 0.000 774.090 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1085.320 4.000 1085.920 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 968.850 1105.025 969.130 1109.025 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 909.970 1105.025 910.250 1109.025 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 427.080 1098.305 427.680 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 201.320 1098.305 201.920 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 595.720 1098.305 596.320 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.090 1105.025 1058.370 1109.025 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 761.850 1105.025 762.130 1109.025 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 193.160 1098.305 193.760 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 507.320 1098.305 507.920 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 91.160 1098.305 91.760 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 771.050 1105.025 771.330 1109.025 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 76.200 1098.305 76.800 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 806.010 1105.025 806.290 1109.025 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 493.720 1098.305 494.320 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 975.160 1098.305 975.760 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.160 4.000 975.760 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1070.360 4.000 1070.960 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.610 1105.025 212.890 1109.025 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 610.680 1098.305 611.280 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 741.240 1098.305 741.840 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1038.770 1105.025 1039.050 1109.025 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 647.770 1105.025 648.050 1109.025 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 608.210 1105.025 608.490 1109.025 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 229.880 1098.305 230.480 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 1105.025 73.970 1109.025 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 682.760 1098.305 683.360 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.450 1105.025 835.730 1109.025 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 624.280 1098.305 624.880 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 858.200 1098.305 858.800 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 747.130 1105.025 747.410 1109.025 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 530.440 1098.305 531.040 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.930 1105.025 485.210 1109.025 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1093.050 1105.025 1093.330 1109.025 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.370 1105.025 54.650 1109.025 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 719.530 0.000 719.810 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 251.640 1098.305 252.240 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 405.810 1105.025 406.090 1109.025 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 791.290 1105.025 791.570 1109.025 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 242.050 1105.025 242.330 1109.025 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 565.800 1098.305 566.400 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.650 1105.025 959.930 1109.025 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 981.730 0.000 982.010 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 722.290 1105.025 722.570 1109.025 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.960 4.000 778.560 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 552.200 1098.305 552.800 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.920 4.000 895.520 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 277.010 1105.025 277.290 1109.025 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 829.640 1098.305 830.240 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.210 1105.025 677.490 1109.025 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 967.010 0.000 967.290 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 840.970 1105.025 841.250 1109.025 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1033.640 1098.305 1034.240 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 187.770 1105.025 188.050 1109.025 ;
    END
  END io_out[9]
  PIN jtag_halt_flag_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1050.730 0.000 1051.010 4.000 ;
    END
  END jtag_halt_flag_i
  PIN jtag_reg_addr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 690.920 1098.305 691.520 ;
    END
  END jtag_reg_addr_i[0]
  PIN jtag_reg_addr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.210 1105.025 148.490 1109.025 ;
    END
  END jtag_reg_addr_i[1]
  PIN jtag_reg_addr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.170 1105.025 390.450 1109.025 ;
    END
  END jtag_reg_addr_i[2]
  PIN jtag_reg_addr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END jtag_reg_addr_i[3]
  PIN jtag_reg_addr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.610 1105.025 143.890 1109.025 ;
    END
  END jtag_reg_addr_i[4]
  PIN jtag_reg_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END jtag_reg_data_i[0]
  PIN jtag_reg_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.930 0.000 784.210 4.000 ;
    END
  END jtag_reg_data_i[10]
  PIN jtag_reg_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 850.170 1105.025 850.450 1109.025 ;
    END
  END jtag_reg_data_i[11]
  PIN jtag_reg_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END jtag_reg_data_i[12]
  PIN jtag_reg_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END jtag_reg_data_i[13]
  PIN jtag_reg_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 939.800 1098.305 940.400 ;
    END
  END jtag_reg_data_i[14]
  PIN jtag_reg_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END jtag_reg_data_i[15]
  PIN jtag_reg_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END jtag_reg_data_i[16]
  PIN jtag_reg_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 578.770 1105.025 579.050 1109.025 ;
    END
  END jtag_reg_data_i[17]
  PIN jtag_reg_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 1105.025 94.210 1109.025 ;
    END
  END jtag_reg_data_i[18]
  PIN jtag_reg_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 449.970 1105.025 450.250 1109.025 ;
    END
  END jtag_reg_data_i[19]
  PIN jtag_reg_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 425.130 1105.025 425.410 1109.025 ;
    END
  END jtag_reg_data_i[1]
  PIN jtag_reg_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 54.440 1098.305 55.040 ;
    END
  END jtag_reg_data_i[20]
  PIN jtag_reg_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.650 1105.025 108.930 1109.025 ;
    END
  END jtag_reg_data_i[21]
  PIN jtag_reg_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 848.330 0.000 848.610 4.000 ;
    END
  END jtag_reg_data_i[22]
  PIN jtag_reg_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 398.520 1098.305 399.120 ;
    END
  END jtag_reg_data_i[23]
  PIN jtag_reg_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.610 1105.025 603.890 1109.025 ;
    END
  END jtag_reg_data_i[24]
  PIN jtag_reg_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 617.480 1098.305 618.080 ;
    END
  END jtag_reg_data_i[25]
  PIN jtag_reg_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END jtag_reg_data_i[26]
  PIN jtag_reg_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END jtag_reg_data_i[27]
  PIN jtag_reg_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END jtag_reg_data_i[28]
  PIN jtag_reg_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END jtag_reg_data_i[29]
  PIN jtag_reg_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END jtag_reg_data_i[2]
  PIN jtag_reg_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 776.570 1105.025 776.850 1109.025 ;
    END
  END jtag_reg_data_i[30]
  PIN jtag_reg_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.250 0.000 803.530 4.000 ;
    END
  END jtag_reg_data_i[31]
  PIN jtag_reg_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 836.440 1098.305 837.040 ;
    END
  END jtag_reg_data_i[3]
  PIN jtag_reg_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1006.570 0.000 1006.850 4.000 ;
    END
  END jtag_reg_data_i[4]
  PIN jtag_reg_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 576.010 0.000 576.290 4.000 ;
    END
  END jtag_reg_data_i[5]
  PIN jtag_reg_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END jtag_reg_data_i[6]
  PIN jtag_reg_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 537.240 1098.305 537.840 ;
    END
  END jtag_reg_data_i[7]
  PIN jtag_reg_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.800 4.000 940.400 ;
    END
  END jtag_reg_data_i[8]
  PIN jtag_reg_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 296.520 1098.305 297.120 ;
    END
  END jtag_reg_data_i[9]
  PIN jtag_reg_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.290 1105.025 860.570 1109.025 ;
    END
  END jtag_reg_data_o[0]
  PIN jtag_reg_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.570 1105.025 316.850 1109.025 ;
    END
  END jtag_reg_data_o[10]
  PIN jtag_reg_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1001.050 0.000 1001.330 4.000 ;
    END
  END jtag_reg_data_o[11]
  PIN jtag_reg_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 826.250 1105.025 826.530 1109.025 ;
    END
  END jtag_reg_data_o[12]
  PIN jtag_reg_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END jtag_reg_data_o[13]
  PIN jtag_reg_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END jtag_reg_data_o[14]
  PIN jtag_reg_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 559.000 1098.305 559.600 ;
    END
  END jtag_reg_data_o[15]
  PIN jtag_reg_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 61.240 1098.305 61.840 ;
    END
  END jtag_reg_data_o[16]
  PIN jtag_reg_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END jtag_reg_data_o[17]
  PIN jtag_reg_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 383.560 1098.305 384.160 ;
    END
  END jtag_reg_data_o[18]
  PIN jtag_reg_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 998.280 1098.305 998.880 ;
    END
  END jtag_reg_data_o[19]
  PIN jtag_reg_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.370 1105.025 445.650 1109.025 ;
    END
  END jtag_reg_data_o[1]
  PIN jtag_reg_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 529.090 1105.025 529.370 1109.025 ;
    END
  END jtag_reg_data_o[20]
  PIN jtag_reg_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END jtag_reg_data_o[21]
  PIN jtag_reg_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 340.040 1098.305 340.640 ;
    END
  END jtag_reg_data_o[22]
  PIN jtag_reg_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END jtag_reg_data_o[23]
  PIN jtag_reg_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 460.090 1105.025 460.370 1109.025 ;
    END
  END jtag_reg_data_o[24]
  PIN jtag_reg_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1100.280 1098.305 1100.880 ;
    END
  END jtag_reg_data_o[25]
  PIN jtag_reg_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 961.560 4.000 962.160 ;
    END
  END jtag_reg_data_o[26]
  PIN jtag_reg_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 518.970 1105.025 519.250 1109.025 ;
    END
  END jtag_reg_data_o[27]
  PIN jtag_reg_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 986.330 0.000 986.610 4.000 ;
    END
  END jtag_reg_data_o[28]
  PIN jtag_reg_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1085.320 1098.305 1085.920 ;
    END
  END jtag_reg_data_o[29]
  PIN jtag_reg_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 568.650 1105.025 568.930 1109.025 ;
    END
  END jtag_reg_data_o[2]
  PIN jtag_reg_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END jtag_reg_data_o[30]
  PIN jtag_reg_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END jtag_reg_data_o[31]
  PIN jtag_reg_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 983.320 1098.305 983.920 ;
    END
  END jtag_reg_data_o[3]
  PIN jtag_reg_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END jtag_reg_data_o[4]
  PIN jtag_reg_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 361.800 1098.305 362.400 ;
    END
  END jtag_reg_data_o[5]
  PIN jtag_reg_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.930 1105.025 163.210 1109.025 ;
    END
  END jtag_reg_data_o[6]
  PIN jtag_reg_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END jtag_reg_data_o[7]
  PIN jtag_reg_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 134.680 1098.305 135.280 ;
    END
  END jtag_reg_data_o[8]
  PIN jtag_reg_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 946.600 1098.305 947.200 ;
    END
  END jtag_reg_data_o[9]
  PIN jtag_reg_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END jtag_reg_we_i
  PIN jtag_reset_flag_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 515.480 1098.305 516.080 ;
    END
  END jtag_reset_flag_i
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 544.040 1098.305 544.640 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 851.400 4.000 852.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.090 1105.025 138.370 1109.025 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 916.680 1098.305 917.280 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 892.490 0.000 892.770 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 953.400 1098.305 954.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 1105.025 15.090 1109.025 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 39.480 1098.305 40.080 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.690 1105.025 533.970 1109.025 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 415.010 1105.025 415.290 1109.025 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1092.120 1098.305 1092.720 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.330 1105.025 227.610 1109.025 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 633.050 1105.025 633.330 1109.025 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 737.010 1105.025 737.290 1109.025 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1080.170 0.000 1080.450 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.490 1105.025 133.770 1109.025 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 844.600 4.000 845.200 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 223.080 1098.305 223.680 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 964.250 1105.025 964.530 1109.025 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 489.530 1105.025 489.810 1109.025 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 1105.025 119.050 1109.025 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 684.570 0.000 684.850 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 781.170 1105.025 781.450 1109.025 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.530 1105.025 98.810 1109.025 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.490 1105.025 271.770 1109.025 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 731.490 1105.025 731.770 1109.025 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 996.450 0.000 996.730 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 439.850 1105.025 440.130 1109.025 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 244.840 1098.305 245.440 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 112.920 1098.305 113.520 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 494.130 1105.025 494.410 1109.025 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 474.810 1105.025 475.090 1109.025 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.570 1105.025 454.850 1109.025 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 712.680 1098.305 713.280 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 588.890 1105.025 589.170 1109.025 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 771.160 1098.305 771.760 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1085.690 0.000 1085.970 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 106.120 1098.305 106.720 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 370.850 1105.025 371.130 1109.025 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 899.850 1105.025 900.130 1109.025 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 691.930 1105.025 692.210 1109.025 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.250 1105.025 113.530 1109.025 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1011.880 1098.305 1012.480 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 756.200 4.000 756.800 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.610 1105.025 1063.890 1109.025 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1041.800 1098.305 1042.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 808.770 0.000 809.050 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 801.410 1105.025 801.690 1109.025 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 376.760 1098.305 377.360 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 463.800 1098.305 464.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 810.610 1105.025 810.890 1109.025 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.610 1105.025 350.890 1109.025 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1060.850 0.000 1061.130 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.930 1105.025 232.210 1109.025 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 500.520 1098.305 501.120 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 208.120 1098.305 208.720 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.130 1105.025 356.410 1109.025 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 17.720 1098.305 18.320 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 360.730 1105.025 361.010 1109.025 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1021.290 0.000 1021.570 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 952.290 0.000 952.570 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 325.080 1098.305 325.680 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 564.050 1105.025 564.330 1109.025 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.080 4.000 903.680 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 214.920 1098.305 215.520 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 870.410 1105.025 870.690 1109.025 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 183.170 1105.025 183.450 1109.025 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1003.810 1105.025 1004.090 1109.025 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 639.240 1098.305 639.840 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 702.050 1105.025 702.330 1109.025 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.160 4.000 873.760 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 1105.025 10.490 1109.025 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.650 1105.025 177.930 1109.025 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.770 1105.025 510.050 1109.025 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 1105.025 59.250 1109.025 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 822.840 1098.305 823.440 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1063.560 1098.305 1064.160 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1070.970 0.000 1071.250 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 1105.025 64.770 1109.025 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 390.360 1098.305 390.960 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1082.930 1105.025 1083.210 1109.025 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 127.880 1098.305 128.480 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 909.880 1098.305 910.480 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.800 4.000 1042.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 675.370 0.000 675.650 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 984.490 1105.025 984.770 1109.025 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 968.360 4.000 968.960 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 142.840 1098.305 143.440 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 897.090 0.000 897.370 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 813.370 0.000 813.650 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 855.690 1105.025 855.970 1109.025 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 669.160 1098.305 669.760 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.410 0.000 1031.690 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.530 1105.025 29.810 1109.025 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 866.360 1098.305 866.960 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 262.290 1105.025 262.570 1109.025 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 164.600 1098.305 165.200 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 429.730 1105.025 430.010 1109.025 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.080 4.000 1005.680 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 553.930 1105.025 554.210 1109.025 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 1105.025 19.690 1109.025 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 97.960 1098.305 98.560 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 875.010 1105.025 875.290 1109.025 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 84.360 1098.305 84.960 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 697.450 1105.025 697.730 1109.025 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.200 4.000 858.800 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 705.880 1098.305 706.480 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 749.400 1098.305 750.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 368.600 1098.305 369.200 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 993.690 1105.025 993.970 1109.025 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 186.360 1098.305 186.960 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 47.640 1098.305 48.240 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 413.480 1098.305 414.080 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 949.530 1105.025 949.810 1109.025 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 266.600 1098.305 267.200 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 954.130 1105.025 954.410 1109.025 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 990.120 1098.305 990.720 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 514.370 1105.025 514.650 1109.025 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 953.400 4.000 954.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.570 1105.025 845.850 1109.025 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1033.250 1105.025 1033.530 1109.025 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1036.010 0.000 1036.290 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 795.890 1105.025 796.170 1109.025 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1026.840 1098.305 1027.440 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 1105.025 25.210 1109.025 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 842.810 0.000 843.090 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 588.920 1098.305 589.520 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 956.890 0.000 957.170 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 173.050 1105.025 173.330 1109.025 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 851.400 1098.305 852.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1040.610 0.000 1040.890 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1068.210 1105.025 1068.490 1109.025 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.130 1105.025 34.410 1109.025 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 301.850 1105.025 302.130 1109.025 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 156.440 1098.305 157.040 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 976.210 0.000 976.490 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 410.410 1105.025 410.690 1109.025 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 318.280 1098.305 318.880 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 887.890 0.000 888.170 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 610.970 0.000 611.250 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 756.330 1105.025 756.610 1109.025 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 687.330 1105.025 687.610 1109.025 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 598.090 1105.025 598.370 1109.025 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 385.570 1105.025 385.850 1109.025 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.170 1105.025 252.450 1109.025 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 331.880 1098.305 332.480 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 471.960 1098.305 472.560 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 777.960 1098.305 778.560 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 346.840 1098.305 347.440 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 549.330 1105.025 549.610 1109.025 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 917.330 0.000 917.610 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 288.360 1098.305 288.960 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1018.530 1105.025 1018.810 1109.025 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1078.330 1105.025 1078.610 1109.025 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.530 1105.025 880.810 1109.025 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 844.600 1098.305 845.200 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 238.040 1098.305 238.640 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 654.200 1098.305 654.800 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 961.560 1098.305 962.160 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 464.690 1105.025 464.970 1109.025 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.010 1105.025 208.290 1109.025 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 741.610 1105.025 741.890 1109.025 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 469.290 1105.025 469.570 1109.025 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.970 1105.025 979.250 1109.025 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 10.920 1098.305 11.520 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 756.200 1098.305 756.800 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.290 1105.025 331.570 1109.025 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.730 1105.025 292.010 1109.025 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.330 1105.025 89.610 1109.025 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.410 1105.025 479.690 1109.025 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1005.080 1098.305 1005.680 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 792.920 1098.305 793.520 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 504.250 1105.025 504.530 1109.025 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 766.450 1105.025 766.730 1109.025 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1013.930 1105.025 1014.210 1109.025 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 281.560 1098.305 282.160 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 499.650 1105.025 499.930 1109.025 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.610 0.000 971.890 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.530 1105.025 1087.810 1109.025 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 1105.025 50.050 1109.025 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 420.280 1098.305 420.880 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 647.400 1098.305 648.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 921.930 0.000 922.210 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 375.450 1105.025 375.730 1109.025 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.610 0.000 902.890 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 914.570 1105.025 914.850 1109.025 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.730 1105.025 223.010 1109.025 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 881.320 1098.305 881.920 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 748.970 0.000 749.250 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1048.600 1098.305 1049.200 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 877.770 0.000 878.050 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 558.530 1105.025 558.810 1109.025 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 920.090 1105.025 920.370 1109.025 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 478.760 1098.305 479.360 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 583.370 1105.025 583.650 1109.025 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1028.650 1105.025 1028.930 1109.025 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 628.450 1105.025 628.730 1109.025 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 734.440 1098.305 735.040 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.890 0.000 1026.170 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.090 1105.025 989.370 1109.025 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 697.720 1098.305 698.320 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.050 1105.025 311.330 1109.025 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1048.600 4.000 1049.200 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.730 0.000 913.010 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 310.120 1098.305 310.720 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 974.370 1105.025 974.650 1109.025 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 820.730 1105.025 821.010 1109.025 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 303.320 1098.305 303.920 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1008.410 1105.025 1008.690 1109.025 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 1105.025 4.970 1109.025 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.810 1105.025 84.090 1109.025 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.130 0.000 655.410 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 682.730 1105.025 683.010 1109.025 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 266.890 1105.025 267.170 1109.025 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 727.640 1098.305 728.240 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 602.520 1098.305 603.120 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 873.160 1098.305 873.760 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.490 1105.025 662.770 1109.025 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 435.250 1105.025 435.530 1109.025 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.370 1105.025 1043.650 1109.025 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 259.800 1098.305 260.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 273.400 1098.305 274.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 637.650 1105.025 637.930 1109.025 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 961.490 0.000 961.770 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 178.200 1098.305 178.800 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 400.290 1105.025 400.570 1109.025 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1047.970 1105.025 1048.250 1109.025 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 895.250 1105.025 895.530 1109.025 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 807.880 1098.305 808.480 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.890 1105.025 336.170 1109.025 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 939.410 1105.025 939.690 1109.025 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.210 0.000 769.490 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.770 1105.025 257.050 1109.025 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.890 1105.025 129.170 1109.025 ;
    END
  END la_oen[9]
  PIN rib_ex_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 643.170 1105.025 643.450 1109.025 ;
    END
  END rib_ex_addr_o[0]
  PIN rib_ex_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 632.440 1098.305 633.040 ;
    END
  END rib_ex_addr_o[10]
  PIN rib_ex_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END rib_ex_addr_o[11]
  PIN rib_ex_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END rib_ex_addr_o[12]
  PIN rib_ex_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 786.120 1098.305 786.720 ;
    END
  END rib_ex_addr_o[13]
  PIN rib_ex_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 751.730 1105.025 752.010 1109.025 ;
    END
  END rib_ex_addr_o[14]
  PIN rib_ex_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 865.810 1105.025 866.090 1109.025 ;
    END
  END rib_ex_addr_o[15]
  PIN rib_ex_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END rib_ex_addr_o[16]
  PIN rib_ex_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 998.280 4.000 998.880 ;
    END
  END rib_ex_addr_o[17]
  PIN rib_ex_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END rib_ex_addr_o[18]
  PIN rib_ex_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END rib_ex_addr_o[19]
  PIN rib_ex_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END rib_ex_addr_o[1]
  PIN rib_ex_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 380.970 1105.025 381.250 1109.025 ;
    END
  END rib_ex_addr_o[20]
  PIN rib_ex_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 816.130 1105.025 816.410 1109.025 ;
    END
  END rib_ex_addr_o[21]
  PIN rib_ex_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.120 4.000 990.720 ;
    END
  END rib_ex_addr_o[22]
  PIN rib_ex_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.690 1105.025 395.970 1109.025 ;
    END
  END rib_ex_addr_o[23]
  PIN rib_ex_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 457.000 1098.305 457.600 ;
    END
  END rib_ex_addr_o[24]
  PIN rib_ex_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 885.130 1105.025 885.410 1109.025 ;
    END
  END rib_ex_addr_o[25]
  PIN rib_ex_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END rib_ex_addr_o[26]
  PIN rib_ex_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END rib_ex_addr_o[27]
  PIN rib_ex_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 618.330 1105.025 618.610 1109.025 ;
    END
  END rib_ex_addr_o[28]
  PIN rib_ex_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 830.850 1105.025 831.130 1109.025 ;
    END
  END rib_ex_addr_o[29]
  PIN rib_ex_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 894.920 1098.305 895.520 ;
    END
  END rib_ex_addr_o[2]
  PIN rib_ex_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1070.360 1098.305 1070.960 ;
    END
  END rib_ex_addr_o[30]
  PIN rib_ex_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 716.770 1105.025 717.050 1109.025 ;
    END
  END rib_ex_addr_o[31]
  PIN rib_ex_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END rib_ex_addr_o[3]
  PIN rib_ex_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END rib_ex_addr_o[4]
  PIN rib_ex_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 539.210 1105.025 539.490 1109.025 ;
    END
  END rib_ex_addr_o[5]
  PIN rib_ex_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END rib_ex_addr_o[6]
  PIN rib_ex_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 946.600 4.000 947.200 ;
    END
  END rib_ex_addr_o[7]
  PIN rib_ex_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END rib_ex_addr_o[8]
  PIN rib_ex_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END rib_ex_addr_o[9]
  PIN rib_ex_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 69.400 1098.305 70.000 ;
    END
  END rib_ex_data_i[0]
  PIN rib_ex_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.760 4.000 1057.360 ;
    END
  END rib_ex_data_i[10]
  PIN rib_ex_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1063.560 4.000 1064.160 ;
    END
  END rib_ex_data_i[11]
  PIN rib_ex_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END rib_ex_data_i[12]
  PIN rib_ex_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 119.720 1098.305 120.320 ;
    END
  END rib_ex_data_i[13]
  PIN rib_ex_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END rib_ex_data_i[14]
  PIN rib_ex_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END rib_ex_data_i[15]
  PIN rib_ex_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.330 0.000 1055.610 4.000 ;
    END
  END rib_ex_data_i[16]
  PIN rib_ex_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.490 0.000 823.770 4.000 ;
    END
  END rib_ex_data_i[17]
  PIN rib_ex_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END rib_ex_data_i[18]
  PIN rib_ex_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END rib_ex_data_i[19]
  PIN rib_ex_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1056.760 1098.305 1057.360 ;
    END
  END rib_ex_data_i[1]
  PIN rib_ex_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 1105.025 39.930 1109.025 ;
    END
  END rib_ex_data_i[20]
  PIN rib_ex_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END rib_ex_data_i[21]
  PIN rib_ex_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END rib_ex_data_i[22]
  PIN rib_ex_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1078.520 1098.305 1079.120 ;
    END
  END rib_ex_data_i[23]
  PIN rib_ex_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END rib_ex_data_i[24]
  PIN rib_ex_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END rib_ex_data_i[25]
  PIN rib_ex_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 778.410 0.000 778.690 4.000 ;
    END
  END rib_ex_data_i[26]
  PIN rib_ex_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END rib_ex_data_i[27]
  PIN rib_ex_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 968.360 1098.305 968.960 ;
    END
  END rib_ex_data_i[28]
  PIN rib_ex_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 622.930 1105.025 623.210 1109.025 ;
    END
  END rib_ex_data_i[29]
  PIN rib_ex_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.210 1105.025 217.490 1109.025 ;
    END
  END rib_ex_data_i[2]
  PIN rib_ex_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 580.760 1098.305 581.360 ;
    END
  END rib_ex_data_i[30]
  PIN rib_ex_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 326.690 1105.025 326.970 1109.025 ;
    END
  END rib_ex_data_i[31]
  PIN rib_ex_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.450 1105.025 237.730 1109.025 ;
    END
  END rib_ex_data_i[3]
  PIN rib_ex_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 612.810 1105.025 613.090 1109.025 ;
    END
  END rib_ex_data_i[4]
  PIN rib_ex_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 306.450 1105.025 306.730 1109.025 ;
    END
  END rib_ex_data_i[5]
  PIN rib_ex_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 661.000 1098.305 661.600 ;
    END
  END rib_ex_data_i[6]
  PIN rib_ex_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END rib_ex_data_i[7]
  PIN rib_ex_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END rib_ex_data_i[8]
  PIN rib_ex_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 828.090 0.000 828.370 4.000 ;
    END
  END rib_ex_data_i[9]
  PIN rib_ex_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 524.490 1105.025 524.770 1109.025 ;
    END
  END rib_ex_data_o[0]
  PIN rib_ex_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END rib_ex_data_o[10]
  PIN rib_ex_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1090.290 0.000 1090.570 4.000 ;
    END
  END rib_ex_data_o[11]
  PIN rib_ex_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 355.000 1098.305 355.600 ;
    END
  END rib_ex_data_o[12]
  PIN rib_ex_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 435.240 1098.305 435.840 ;
    END
  END rib_ex_data_o[13]
  PIN rib_ex_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 485.560 1098.305 486.160 ;
    END
  END rib_ex_data_o[14]
  PIN rib_ex_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.330 1105.025 296.610 1109.025 ;
    END
  END rib_ex_data_o[15]
  PIN rib_ex_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1092.120 4.000 1092.720 ;
    END
  END rib_ex_data_o[16]
  PIN rib_ex_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 905.370 1105.025 905.650 1109.025 ;
    END
  END rib_ex_data_o[17]
  PIN rib_ex_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END rib_ex_data_o[18]
  PIN rib_ex_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 675.960 1098.305 676.560 ;
    END
  END rib_ex_data_o[19]
  PIN rib_ex_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END rib_ex_data_o[1]
  PIN rib_ex_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END rib_ex_data_o[20]
  PIN rib_ex_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 192.370 1105.025 192.650 1109.025 ;
    END
  END rib_ex_data_o[21]
  PIN rib_ex_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 707.570 1105.025 707.850 1109.025 ;
    END
  END rib_ex_data_o[22]
  PIN rib_ex_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END rib_ex_data_o[23]
  PIN rib_ex_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.690 1105.025 924.970 1109.025 ;
    END
  END rib_ex_data_o[24]
  PIN rib_ex_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END rib_ex_data_o[25]
  PIN rib_ex_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END rib_ex_data_o[26]
  PIN rib_ex_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.410 1105.025 341.690 1109.025 ;
    END
  END rib_ex_data_o[27]
  PIN rib_ex_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 903.080 1098.305 903.680 ;
    END
  END rib_ex_data_o[28]
  PIN rib_ex_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END rib_ex_data_o[29]
  PIN rib_ex_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 764.360 1098.305 764.960 ;
    END
  END rib_ex_data_o[2]
  PIN rib_ex_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.450 1105.025 168.730 1109.025 ;
    END
  END rib_ex_data_o[30]
  PIN rib_ex_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END rib_ex_data_o[31]
  PIN rib_ex_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END rib_ex_data_o[3]
  PIN rib_ex_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 719.480 1098.305 720.080 ;
    END
  END rib_ex_data_o[4]
  PIN rib_ex_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END rib_ex_data_o[5]
  PIN rib_ex_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 652.370 1105.025 652.650 1109.025 ;
    END
  END rib_ex_data_o[6]
  PIN rib_ex_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END rib_ex_data_o[7]
  PIN rib_ex_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END rib_ex_data_o[8]
  PIN rib_ex_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END rib_ex_data_o[9]
  PIN rib_ex_req_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END rib_ex_req_o
  PIN rib_ex_we_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.170 1105.025 321.450 1109.025 ;
    END
  END rib_ex_we_o
  PIN rib_hold_flag_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 833.610 0.000 833.890 4.000 ;
    END
  END rib_hold_flag_i
  PIN rib_pc_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1065.450 0.000 1065.730 4.000 ;
    END
  END rib_pc_addr_o[0]
  PIN rib_pc_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.050 1105.025 1024.330 1109.025 ;
    END
  END rib_pc_addr_o[10]
  PIN rib_pc_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 442.040 1098.305 442.640 ;
    END
  END rib_pc_addr_o[11]
  PIN rib_pc_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 694.690 0.000 694.970 4.000 ;
    END
  END rib_pc_addr_o[12]
  PIN rib_pc_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 448.840 1098.305 449.440 ;
    END
  END rib_pc_addr_o[13]
  PIN rib_pc_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.160 4.000 771.760 ;
    END
  END rib_pc_addr_o[14]
  PIN rib_pc_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.810 1105.025 153.090 1109.025 ;
    END
  END rib_pc_addr_o[15]
  PIN rib_pc_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 522.280 1098.305 522.880 ;
    END
  END rib_pc_addr_o[16]
  PIN rib_pc_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 931.640 1098.305 932.240 ;
    END
  END rib_pc_addr_o[17]
  PIN rib_pc_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 659.730 0.000 660.010 4.000 ;
    END
  END rib_pc_addr_o[18]
  PIN rib_pc_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END rib_pc_addr_o[19]
  PIN rib_pc_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END rib_pc_addr_o[1]
  PIN rib_pc_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.130 1105.025 287.410 1109.025 ;
    END
  END rib_pc_addr_o[20]
  PIN rib_pc_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END rib_pc_addr_o[21]
  PIN rib_pc_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 814.680 1098.305 815.280 ;
    END
  END rib_pc_addr_o[22]
  PIN rib_pc_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 4.000 ;
    END
  END rib_pc_addr_o[23]
  PIN rib_pc_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END rib_pc_addr_o[24]
  PIN rib_pc_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 657.890 1105.025 658.170 1109.025 ;
    END
  END rib_pc_addr_o[25]
  PIN rib_pc_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1100.280 4.000 1100.880 ;
    END
  END rib_pc_addr_o[26]
  PIN rib_pc_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 889.730 1105.025 890.010 1109.025 ;
    END
  END rib_pc_addr_o[27]
  PIN rib_pc_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 1105.025 69.370 1109.025 ;
    END
  END rib_pc_addr_o[28]
  PIN rib_pc_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1094.305 1020.040 1098.305 1020.640 ;
    END
  END rib_pc_addr_o[29]
  PIN rib_pc_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 1105.025 104.330 1109.025 ;
    END
  END rib_pc_addr_o[2]
  PIN rib_pc_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END rib_pc_addr_o[30]
  PIN rib_pc_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END rib_pc_addr_o[31]
  PIN rib_pc_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.690 1105.025 786.970 1109.025 ;
    END
  END rib_pc_addr_o[3]
  PIN rib_pc_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 4.000 917.280 ;
    END
  END rib_pc_addr_o[4]
  PIN rib_pc_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1072.810 1105.025 1073.090 1109.025 ;
    END
  END rib_pc_addr_o[5]
  PIN rib_pc_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 346.010 1105.025 346.290 1109.025 ;
    END
  END rib_pc_addr_o[6]
  PIN rib_pc_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 999.210 1105.025 999.490 1109.025 ;
    END
  END rib_pc_addr_o[7]
  PIN rib_pc_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 366.250 1105.025 366.530 1109.025 ;
    END
  END rib_pc_addr_o[8]
  PIN rib_pc_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 247.570 1105.025 247.850 1109.025 ;
    END
  END rib_pc_addr_o[9]
  PIN rib_pc_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END rib_pc_data_i[0]
  PIN rib_pc_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 171.400 1098.305 172.000 ;
    END
  END rib_pc_data_i[10]
  PIN rib_pc_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.890 1105.025 198.170 1109.025 ;
    END
  END rib_pc_data_i[11]
  PIN rib_pc_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END rib_pc_data_i[12]
  PIN rib_pc_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END rib_pc_data_i[13]
  PIN rib_pc_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 799.720 1098.305 800.320 ;
    END
  END rib_pc_data_i[14]
  PIN rib_pc_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1078.520 4.000 1079.120 ;
    END
  END rib_pc_data_i[15]
  PIN rib_pc_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 888.120 1098.305 888.720 ;
    END
  END rib_pc_data_i[16]
  PIN rib_pc_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END rib_pc_data_i[17]
  PIN rib_pc_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.530 1105.025 420.810 1109.025 ;
    END
  END rib_pc_data_i[18]
  PIN rib_pc_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 25.880 1098.305 26.480 ;
    END
  END rib_pc_data_i[19]
  PIN rib_pc_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 573.250 1105.025 573.530 1109.025 ;
    END
  END rib_pc_data_i[1]
  PIN rib_pc_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 873.170 0.000 873.450 4.000 ;
    END
  END rib_pc_data_i[20]
  PIN rib_pc_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END rib_pc_data_i[21]
  PIN rib_pc_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END rib_pc_data_i[22]
  PIN rib_pc_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 764.360 4.000 764.960 ;
    END
  END rib_pc_data_i[23]
  PIN rib_pc_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END rib_pc_data_i[24]
  PIN rib_pc_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 1105.025 79.490 1109.025 ;
    END
  END rib_pc_data_i[25]
  PIN rib_pc_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.010 1105.025 668.290 1109.025 ;
    END
  END rib_pc_data_i[26]
  PIN rib_pc_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 573.960 1098.305 574.560 ;
    END
  END rib_pc_data_i[27]
  PIN rib_pc_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END rib_pc_data_i[28]
  PIN rib_pc_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END rib_pc_data_i[29]
  PIN rib_pc_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 712.170 1105.025 712.450 1109.025 ;
    END
  END rib_pc_data_i[2]
  PIN rib_pc_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.290 1105.025 929.570 1109.025 ;
    END
  END rib_pc_data_i[30]
  PIN rib_pc_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1053.490 1105.025 1053.770 1109.025 ;
    END
  END rib_pc_data_i[31]
  PIN rib_pc_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.330 1105.025 158.610 1109.025 ;
    END
  END rib_pc_data_i[3]
  PIN rib_pc_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END rib_pc_data_i[4]
  PIN rib_pc_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 944.930 1105.025 945.210 1109.025 ;
    END
  END rib_pc_data_i[5]
  PIN rib_pc_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END rib_pc_data_i[6]
  PIN rib_pc_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1094.305 149.640 1098.305 150.240 ;
    END
  END rib_pc_data_i[7]
  PIN rib_pc_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END rib_pc_data_i[8]
  PIN rib_pc_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 726.890 1105.025 727.170 1109.025 ;
    END
  END rib_pc_data_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 593.490 1105.025 593.770 1109.025 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 4.000 ;
    END
  END wb_rst_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 1092.500 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 1092.500 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1092.500 1096.245 ;
      LAYER met1 ;
        RECT 2.830 5.820 1093.350 1097.480 ;
      LAYER met2 ;
        RECT 2.860 1104.745 4.410 1105.025 ;
        RECT 5.250 1104.745 9.930 1105.025 ;
        RECT 10.770 1104.745 14.530 1105.025 ;
        RECT 15.370 1104.745 19.130 1105.025 ;
        RECT 19.970 1104.745 24.650 1105.025 ;
        RECT 25.490 1104.745 29.250 1105.025 ;
        RECT 30.090 1104.745 33.850 1105.025 ;
        RECT 34.690 1104.745 39.370 1105.025 ;
        RECT 40.210 1104.745 43.970 1105.025 ;
        RECT 44.810 1104.745 49.490 1105.025 ;
        RECT 50.330 1104.745 54.090 1105.025 ;
        RECT 54.930 1104.745 58.690 1105.025 ;
        RECT 59.530 1104.745 64.210 1105.025 ;
        RECT 65.050 1104.745 68.810 1105.025 ;
        RECT 69.650 1104.745 73.410 1105.025 ;
        RECT 74.250 1104.745 78.930 1105.025 ;
        RECT 79.770 1104.745 83.530 1105.025 ;
        RECT 84.370 1104.745 89.050 1105.025 ;
        RECT 89.890 1104.745 93.650 1105.025 ;
        RECT 94.490 1104.745 98.250 1105.025 ;
        RECT 99.090 1104.745 103.770 1105.025 ;
        RECT 104.610 1104.745 108.370 1105.025 ;
        RECT 109.210 1104.745 112.970 1105.025 ;
        RECT 113.810 1104.745 118.490 1105.025 ;
        RECT 119.330 1104.745 123.090 1105.025 ;
        RECT 123.930 1104.745 128.610 1105.025 ;
        RECT 129.450 1104.745 133.210 1105.025 ;
        RECT 134.050 1104.745 137.810 1105.025 ;
        RECT 138.650 1104.745 143.330 1105.025 ;
        RECT 144.170 1104.745 147.930 1105.025 ;
        RECT 148.770 1104.745 152.530 1105.025 ;
        RECT 153.370 1104.745 158.050 1105.025 ;
        RECT 158.890 1104.745 162.650 1105.025 ;
        RECT 163.490 1104.745 168.170 1105.025 ;
        RECT 169.010 1104.745 172.770 1105.025 ;
        RECT 173.610 1104.745 177.370 1105.025 ;
        RECT 178.210 1104.745 182.890 1105.025 ;
        RECT 183.730 1104.745 187.490 1105.025 ;
        RECT 188.330 1104.745 192.090 1105.025 ;
        RECT 192.930 1104.745 197.610 1105.025 ;
        RECT 198.450 1104.745 202.210 1105.025 ;
        RECT 203.050 1104.745 207.730 1105.025 ;
        RECT 208.570 1104.745 212.330 1105.025 ;
        RECT 213.170 1104.745 216.930 1105.025 ;
        RECT 217.770 1104.745 222.450 1105.025 ;
        RECT 223.290 1104.745 227.050 1105.025 ;
        RECT 227.890 1104.745 231.650 1105.025 ;
        RECT 232.490 1104.745 237.170 1105.025 ;
        RECT 238.010 1104.745 241.770 1105.025 ;
        RECT 242.610 1104.745 247.290 1105.025 ;
        RECT 248.130 1104.745 251.890 1105.025 ;
        RECT 252.730 1104.745 256.490 1105.025 ;
        RECT 257.330 1104.745 262.010 1105.025 ;
        RECT 262.850 1104.745 266.610 1105.025 ;
        RECT 267.450 1104.745 271.210 1105.025 ;
        RECT 272.050 1104.745 276.730 1105.025 ;
        RECT 277.570 1104.745 281.330 1105.025 ;
        RECT 282.170 1104.745 286.850 1105.025 ;
        RECT 287.690 1104.745 291.450 1105.025 ;
        RECT 292.290 1104.745 296.050 1105.025 ;
        RECT 296.890 1104.745 301.570 1105.025 ;
        RECT 302.410 1104.745 306.170 1105.025 ;
        RECT 307.010 1104.745 310.770 1105.025 ;
        RECT 311.610 1104.745 316.290 1105.025 ;
        RECT 317.130 1104.745 320.890 1105.025 ;
        RECT 321.730 1104.745 326.410 1105.025 ;
        RECT 327.250 1104.745 331.010 1105.025 ;
        RECT 331.850 1104.745 335.610 1105.025 ;
        RECT 336.450 1104.745 341.130 1105.025 ;
        RECT 341.970 1104.745 345.730 1105.025 ;
        RECT 346.570 1104.745 350.330 1105.025 ;
        RECT 351.170 1104.745 355.850 1105.025 ;
        RECT 356.690 1104.745 360.450 1105.025 ;
        RECT 361.290 1104.745 365.970 1105.025 ;
        RECT 366.810 1104.745 370.570 1105.025 ;
        RECT 371.410 1104.745 375.170 1105.025 ;
        RECT 376.010 1104.745 380.690 1105.025 ;
        RECT 381.530 1104.745 385.290 1105.025 ;
        RECT 386.130 1104.745 389.890 1105.025 ;
        RECT 390.730 1104.745 395.410 1105.025 ;
        RECT 396.250 1104.745 400.010 1105.025 ;
        RECT 400.850 1104.745 405.530 1105.025 ;
        RECT 406.370 1104.745 410.130 1105.025 ;
        RECT 410.970 1104.745 414.730 1105.025 ;
        RECT 415.570 1104.745 420.250 1105.025 ;
        RECT 421.090 1104.745 424.850 1105.025 ;
        RECT 425.690 1104.745 429.450 1105.025 ;
        RECT 430.290 1104.745 434.970 1105.025 ;
        RECT 435.810 1104.745 439.570 1105.025 ;
        RECT 440.410 1104.745 445.090 1105.025 ;
        RECT 445.930 1104.745 449.690 1105.025 ;
        RECT 450.530 1104.745 454.290 1105.025 ;
        RECT 455.130 1104.745 459.810 1105.025 ;
        RECT 460.650 1104.745 464.410 1105.025 ;
        RECT 465.250 1104.745 469.010 1105.025 ;
        RECT 469.850 1104.745 474.530 1105.025 ;
        RECT 475.370 1104.745 479.130 1105.025 ;
        RECT 479.970 1104.745 484.650 1105.025 ;
        RECT 485.490 1104.745 489.250 1105.025 ;
        RECT 490.090 1104.745 493.850 1105.025 ;
        RECT 494.690 1104.745 499.370 1105.025 ;
        RECT 500.210 1104.745 503.970 1105.025 ;
        RECT 504.810 1104.745 509.490 1105.025 ;
        RECT 510.330 1104.745 514.090 1105.025 ;
        RECT 514.930 1104.745 518.690 1105.025 ;
        RECT 519.530 1104.745 524.210 1105.025 ;
        RECT 525.050 1104.745 528.810 1105.025 ;
        RECT 529.650 1104.745 533.410 1105.025 ;
        RECT 534.250 1104.745 538.930 1105.025 ;
        RECT 539.770 1104.745 543.530 1105.025 ;
        RECT 544.370 1104.745 549.050 1105.025 ;
        RECT 549.890 1104.745 553.650 1105.025 ;
        RECT 554.490 1104.745 558.250 1105.025 ;
        RECT 559.090 1104.745 563.770 1105.025 ;
        RECT 564.610 1104.745 568.370 1105.025 ;
        RECT 569.210 1104.745 572.970 1105.025 ;
        RECT 573.810 1104.745 578.490 1105.025 ;
        RECT 579.330 1104.745 583.090 1105.025 ;
        RECT 583.930 1104.745 588.610 1105.025 ;
        RECT 589.450 1104.745 593.210 1105.025 ;
        RECT 594.050 1104.745 597.810 1105.025 ;
        RECT 598.650 1104.745 603.330 1105.025 ;
        RECT 604.170 1104.745 607.930 1105.025 ;
        RECT 608.770 1104.745 612.530 1105.025 ;
        RECT 613.370 1104.745 618.050 1105.025 ;
        RECT 618.890 1104.745 622.650 1105.025 ;
        RECT 623.490 1104.745 628.170 1105.025 ;
        RECT 629.010 1104.745 632.770 1105.025 ;
        RECT 633.610 1104.745 637.370 1105.025 ;
        RECT 638.210 1104.745 642.890 1105.025 ;
        RECT 643.730 1104.745 647.490 1105.025 ;
        RECT 648.330 1104.745 652.090 1105.025 ;
        RECT 652.930 1104.745 657.610 1105.025 ;
        RECT 658.450 1104.745 662.210 1105.025 ;
        RECT 663.050 1104.745 667.730 1105.025 ;
        RECT 668.570 1104.745 672.330 1105.025 ;
        RECT 673.170 1104.745 676.930 1105.025 ;
        RECT 677.770 1104.745 682.450 1105.025 ;
        RECT 683.290 1104.745 687.050 1105.025 ;
        RECT 687.890 1104.745 691.650 1105.025 ;
        RECT 692.490 1104.745 697.170 1105.025 ;
        RECT 698.010 1104.745 701.770 1105.025 ;
        RECT 702.610 1104.745 707.290 1105.025 ;
        RECT 708.130 1104.745 711.890 1105.025 ;
        RECT 712.730 1104.745 716.490 1105.025 ;
        RECT 717.330 1104.745 722.010 1105.025 ;
        RECT 722.850 1104.745 726.610 1105.025 ;
        RECT 727.450 1104.745 731.210 1105.025 ;
        RECT 732.050 1104.745 736.730 1105.025 ;
        RECT 737.570 1104.745 741.330 1105.025 ;
        RECT 742.170 1104.745 746.850 1105.025 ;
        RECT 747.690 1104.745 751.450 1105.025 ;
        RECT 752.290 1104.745 756.050 1105.025 ;
        RECT 756.890 1104.745 761.570 1105.025 ;
        RECT 762.410 1104.745 766.170 1105.025 ;
        RECT 767.010 1104.745 770.770 1105.025 ;
        RECT 771.610 1104.745 776.290 1105.025 ;
        RECT 777.130 1104.745 780.890 1105.025 ;
        RECT 781.730 1104.745 786.410 1105.025 ;
        RECT 787.250 1104.745 791.010 1105.025 ;
        RECT 791.850 1104.745 795.610 1105.025 ;
        RECT 796.450 1104.745 801.130 1105.025 ;
        RECT 801.970 1104.745 805.730 1105.025 ;
        RECT 806.570 1104.745 810.330 1105.025 ;
        RECT 811.170 1104.745 815.850 1105.025 ;
        RECT 816.690 1104.745 820.450 1105.025 ;
        RECT 821.290 1104.745 825.970 1105.025 ;
        RECT 826.810 1104.745 830.570 1105.025 ;
        RECT 831.410 1104.745 835.170 1105.025 ;
        RECT 836.010 1104.745 840.690 1105.025 ;
        RECT 841.530 1104.745 845.290 1105.025 ;
        RECT 846.130 1104.745 849.890 1105.025 ;
        RECT 850.730 1104.745 855.410 1105.025 ;
        RECT 856.250 1104.745 860.010 1105.025 ;
        RECT 860.850 1104.745 865.530 1105.025 ;
        RECT 866.370 1104.745 870.130 1105.025 ;
        RECT 870.970 1104.745 874.730 1105.025 ;
        RECT 875.570 1104.745 880.250 1105.025 ;
        RECT 881.090 1104.745 884.850 1105.025 ;
        RECT 885.690 1104.745 889.450 1105.025 ;
        RECT 890.290 1104.745 894.970 1105.025 ;
        RECT 895.810 1104.745 899.570 1105.025 ;
        RECT 900.410 1104.745 905.090 1105.025 ;
        RECT 905.930 1104.745 909.690 1105.025 ;
        RECT 910.530 1104.745 914.290 1105.025 ;
        RECT 915.130 1104.745 919.810 1105.025 ;
        RECT 920.650 1104.745 924.410 1105.025 ;
        RECT 925.250 1104.745 929.010 1105.025 ;
        RECT 929.850 1104.745 934.530 1105.025 ;
        RECT 935.370 1104.745 939.130 1105.025 ;
        RECT 939.970 1104.745 944.650 1105.025 ;
        RECT 945.490 1104.745 949.250 1105.025 ;
        RECT 950.090 1104.745 953.850 1105.025 ;
        RECT 954.690 1104.745 959.370 1105.025 ;
        RECT 960.210 1104.745 963.970 1105.025 ;
        RECT 964.810 1104.745 968.570 1105.025 ;
        RECT 969.410 1104.745 974.090 1105.025 ;
        RECT 974.930 1104.745 978.690 1105.025 ;
        RECT 979.530 1104.745 984.210 1105.025 ;
        RECT 985.050 1104.745 988.810 1105.025 ;
        RECT 989.650 1104.745 993.410 1105.025 ;
        RECT 994.250 1104.745 998.930 1105.025 ;
        RECT 999.770 1104.745 1003.530 1105.025 ;
        RECT 1004.370 1104.745 1008.130 1105.025 ;
        RECT 1008.970 1104.745 1013.650 1105.025 ;
        RECT 1014.490 1104.745 1018.250 1105.025 ;
        RECT 1019.090 1104.745 1023.770 1105.025 ;
        RECT 1024.610 1104.745 1028.370 1105.025 ;
        RECT 1029.210 1104.745 1032.970 1105.025 ;
        RECT 1033.810 1104.745 1038.490 1105.025 ;
        RECT 1039.330 1104.745 1043.090 1105.025 ;
        RECT 1043.930 1104.745 1047.690 1105.025 ;
        RECT 1048.530 1104.745 1053.210 1105.025 ;
        RECT 1054.050 1104.745 1057.810 1105.025 ;
        RECT 1058.650 1104.745 1063.330 1105.025 ;
        RECT 1064.170 1104.745 1067.930 1105.025 ;
        RECT 1068.770 1104.745 1072.530 1105.025 ;
        RECT 1073.370 1104.745 1078.050 1105.025 ;
        RECT 1078.890 1104.745 1082.650 1105.025 ;
        RECT 1083.490 1104.745 1087.250 1105.025 ;
        RECT 1088.090 1104.745 1092.770 1105.025 ;
        RECT 2.860 4.280 1093.320 1104.745 ;
        RECT 3.410 4.000 7.170 4.280 ;
        RECT 8.010 4.000 11.770 4.280 ;
        RECT 12.610 4.000 17.290 4.280 ;
        RECT 18.130 4.000 21.890 4.280 ;
        RECT 22.730 4.000 26.490 4.280 ;
        RECT 27.330 4.000 32.010 4.280 ;
        RECT 32.850 4.000 36.610 4.280 ;
        RECT 37.450 4.000 42.130 4.280 ;
        RECT 42.970 4.000 46.730 4.280 ;
        RECT 47.570 4.000 51.330 4.280 ;
        RECT 52.170 4.000 56.850 4.280 ;
        RECT 57.690 4.000 61.450 4.280 ;
        RECT 62.290 4.000 66.050 4.280 ;
        RECT 66.890 4.000 71.570 4.280 ;
        RECT 72.410 4.000 76.170 4.280 ;
        RECT 77.010 4.000 81.690 4.280 ;
        RECT 82.530 4.000 86.290 4.280 ;
        RECT 87.130 4.000 90.890 4.280 ;
        RECT 91.730 4.000 96.410 4.280 ;
        RECT 97.250 4.000 101.010 4.280 ;
        RECT 101.850 4.000 105.610 4.280 ;
        RECT 106.450 4.000 111.130 4.280 ;
        RECT 111.970 4.000 115.730 4.280 ;
        RECT 116.570 4.000 121.250 4.280 ;
        RECT 122.090 4.000 125.850 4.280 ;
        RECT 126.690 4.000 130.450 4.280 ;
        RECT 131.290 4.000 135.970 4.280 ;
        RECT 136.810 4.000 140.570 4.280 ;
        RECT 141.410 4.000 145.170 4.280 ;
        RECT 146.010 4.000 150.690 4.280 ;
        RECT 151.530 4.000 155.290 4.280 ;
        RECT 156.130 4.000 160.810 4.280 ;
        RECT 161.650 4.000 165.410 4.280 ;
        RECT 166.250 4.000 170.010 4.280 ;
        RECT 170.850 4.000 175.530 4.280 ;
        RECT 176.370 4.000 180.130 4.280 ;
        RECT 180.970 4.000 184.730 4.280 ;
        RECT 185.570 4.000 190.250 4.280 ;
        RECT 191.090 4.000 194.850 4.280 ;
        RECT 195.690 4.000 200.370 4.280 ;
        RECT 201.210 4.000 204.970 4.280 ;
        RECT 205.810 4.000 209.570 4.280 ;
        RECT 210.410 4.000 215.090 4.280 ;
        RECT 215.930 4.000 219.690 4.280 ;
        RECT 220.530 4.000 224.290 4.280 ;
        RECT 225.130 4.000 229.810 4.280 ;
        RECT 230.650 4.000 234.410 4.280 ;
        RECT 235.250 4.000 239.930 4.280 ;
        RECT 240.770 4.000 244.530 4.280 ;
        RECT 245.370 4.000 249.130 4.280 ;
        RECT 249.970 4.000 254.650 4.280 ;
        RECT 255.490 4.000 259.250 4.280 ;
        RECT 260.090 4.000 263.850 4.280 ;
        RECT 264.690 4.000 269.370 4.280 ;
        RECT 270.210 4.000 273.970 4.280 ;
        RECT 274.810 4.000 279.490 4.280 ;
        RECT 280.330 4.000 284.090 4.280 ;
        RECT 284.930 4.000 288.690 4.280 ;
        RECT 289.530 4.000 294.210 4.280 ;
        RECT 295.050 4.000 298.810 4.280 ;
        RECT 299.650 4.000 303.410 4.280 ;
        RECT 304.250 4.000 308.930 4.280 ;
        RECT 309.770 4.000 313.530 4.280 ;
        RECT 314.370 4.000 319.050 4.280 ;
        RECT 319.890 4.000 323.650 4.280 ;
        RECT 324.490 4.000 328.250 4.280 ;
        RECT 329.090 4.000 333.770 4.280 ;
        RECT 334.610 4.000 338.370 4.280 ;
        RECT 339.210 4.000 342.970 4.280 ;
        RECT 343.810 4.000 348.490 4.280 ;
        RECT 349.330 4.000 353.090 4.280 ;
        RECT 353.930 4.000 358.610 4.280 ;
        RECT 359.450 4.000 363.210 4.280 ;
        RECT 364.050 4.000 367.810 4.280 ;
        RECT 368.650 4.000 373.330 4.280 ;
        RECT 374.170 4.000 377.930 4.280 ;
        RECT 378.770 4.000 382.530 4.280 ;
        RECT 383.370 4.000 388.050 4.280 ;
        RECT 388.890 4.000 392.650 4.280 ;
        RECT 393.490 4.000 398.170 4.280 ;
        RECT 399.010 4.000 402.770 4.280 ;
        RECT 403.610 4.000 407.370 4.280 ;
        RECT 408.210 4.000 412.890 4.280 ;
        RECT 413.730 4.000 417.490 4.280 ;
        RECT 418.330 4.000 422.090 4.280 ;
        RECT 422.930 4.000 427.610 4.280 ;
        RECT 428.450 4.000 432.210 4.280 ;
        RECT 433.050 4.000 437.730 4.280 ;
        RECT 438.570 4.000 442.330 4.280 ;
        RECT 443.170 4.000 446.930 4.280 ;
        RECT 447.770 4.000 452.450 4.280 ;
        RECT 453.290 4.000 457.050 4.280 ;
        RECT 457.890 4.000 461.650 4.280 ;
        RECT 462.490 4.000 467.170 4.280 ;
        RECT 468.010 4.000 471.770 4.280 ;
        RECT 472.610 4.000 477.290 4.280 ;
        RECT 478.130 4.000 481.890 4.280 ;
        RECT 482.730 4.000 486.490 4.280 ;
        RECT 487.330 4.000 492.010 4.280 ;
        RECT 492.850 4.000 496.610 4.280 ;
        RECT 497.450 4.000 501.210 4.280 ;
        RECT 502.050 4.000 506.730 4.280 ;
        RECT 507.570 4.000 511.330 4.280 ;
        RECT 512.170 4.000 516.850 4.280 ;
        RECT 517.690 4.000 521.450 4.280 ;
        RECT 522.290 4.000 526.050 4.280 ;
        RECT 526.890 4.000 531.570 4.280 ;
        RECT 532.410 4.000 536.170 4.280 ;
        RECT 537.010 4.000 540.770 4.280 ;
        RECT 541.610 4.000 546.290 4.280 ;
        RECT 547.130 4.000 550.890 4.280 ;
        RECT 551.730 4.000 556.410 4.280 ;
        RECT 557.250 4.000 561.010 4.280 ;
        RECT 561.850 4.000 565.610 4.280 ;
        RECT 566.450 4.000 571.130 4.280 ;
        RECT 571.970 4.000 575.730 4.280 ;
        RECT 576.570 4.000 580.330 4.280 ;
        RECT 581.170 4.000 585.850 4.280 ;
        RECT 586.690 4.000 590.450 4.280 ;
        RECT 591.290 4.000 595.970 4.280 ;
        RECT 596.810 4.000 600.570 4.280 ;
        RECT 601.410 4.000 605.170 4.280 ;
        RECT 606.010 4.000 610.690 4.280 ;
        RECT 611.530 4.000 615.290 4.280 ;
        RECT 616.130 4.000 619.890 4.280 ;
        RECT 620.730 4.000 625.410 4.280 ;
        RECT 626.250 4.000 630.010 4.280 ;
        RECT 630.850 4.000 635.530 4.280 ;
        RECT 636.370 4.000 640.130 4.280 ;
        RECT 640.970 4.000 644.730 4.280 ;
        RECT 645.570 4.000 650.250 4.280 ;
        RECT 651.090 4.000 654.850 4.280 ;
        RECT 655.690 4.000 659.450 4.280 ;
        RECT 660.290 4.000 664.970 4.280 ;
        RECT 665.810 4.000 669.570 4.280 ;
        RECT 670.410 4.000 675.090 4.280 ;
        RECT 675.930 4.000 679.690 4.280 ;
        RECT 680.530 4.000 684.290 4.280 ;
        RECT 685.130 4.000 689.810 4.280 ;
        RECT 690.650 4.000 694.410 4.280 ;
        RECT 695.250 4.000 699.010 4.280 ;
        RECT 699.850 4.000 704.530 4.280 ;
        RECT 705.370 4.000 709.130 4.280 ;
        RECT 709.970 4.000 714.650 4.280 ;
        RECT 715.490 4.000 719.250 4.280 ;
        RECT 720.090 4.000 723.850 4.280 ;
        RECT 724.690 4.000 729.370 4.280 ;
        RECT 730.210 4.000 733.970 4.280 ;
        RECT 734.810 4.000 738.570 4.280 ;
        RECT 739.410 4.000 744.090 4.280 ;
        RECT 744.930 4.000 748.690 4.280 ;
        RECT 749.530 4.000 754.210 4.280 ;
        RECT 755.050 4.000 758.810 4.280 ;
        RECT 759.650 4.000 763.410 4.280 ;
        RECT 764.250 4.000 768.930 4.280 ;
        RECT 769.770 4.000 773.530 4.280 ;
        RECT 774.370 4.000 778.130 4.280 ;
        RECT 778.970 4.000 783.650 4.280 ;
        RECT 784.490 4.000 788.250 4.280 ;
        RECT 789.090 4.000 793.770 4.280 ;
        RECT 794.610 4.000 798.370 4.280 ;
        RECT 799.210 4.000 802.970 4.280 ;
        RECT 803.810 4.000 808.490 4.280 ;
        RECT 809.330 4.000 813.090 4.280 ;
        RECT 813.930 4.000 817.690 4.280 ;
        RECT 818.530 4.000 823.210 4.280 ;
        RECT 824.050 4.000 827.810 4.280 ;
        RECT 828.650 4.000 833.330 4.280 ;
        RECT 834.170 4.000 837.930 4.280 ;
        RECT 838.770 4.000 842.530 4.280 ;
        RECT 843.370 4.000 848.050 4.280 ;
        RECT 848.890 4.000 852.650 4.280 ;
        RECT 853.490 4.000 857.250 4.280 ;
        RECT 858.090 4.000 862.770 4.280 ;
        RECT 863.610 4.000 867.370 4.280 ;
        RECT 868.210 4.000 872.890 4.280 ;
        RECT 873.730 4.000 877.490 4.280 ;
        RECT 878.330 4.000 882.090 4.280 ;
        RECT 882.930 4.000 887.610 4.280 ;
        RECT 888.450 4.000 892.210 4.280 ;
        RECT 893.050 4.000 896.810 4.280 ;
        RECT 897.650 4.000 902.330 4.280 ;
        RECT 903.170 4.000 906.930 4.280 ;
        RECT 907.770 4.000 912.450 4.280 ;
        RECT 913.290 4.000 917.050 4.280 ;
        RECT 917.890 4.000 921.650 4.280 ;
        RECT 922.490 4.000 927.170 4.280 ;
        RECT 928.010 4.000 931.770 4.280 ;
        RECT 932.610 4.000 936.370 4.280 ;
        RECT 937.210 4.000 941.890 4.280 ;
        RECT 942.730 4.000 946.490 4.280 ;
        RECT 947.330 4.000 952.010 4.280 ;
        RECT 952.850 4.000 956.610 4.280 ;
        RECT 957.450 4.000 961.210 4.280 ;
        RECT 962.050 4.000 966.730 4.280 ;
        RECT 967.570 4.000 971.330 4.280 ;
        RECT 972.170 4.000 975.930 4.280 ;
        RECT 976.770 4.000 981.450 4.280 ;
        RECT 982.290 4.000 986.050 4.280 ;
        RECT 986.890 4.000 991.570 4.280 ;
        RECT 992.410 4.000 996.170 4.280 ;
        RECT 997.010 4.000 1000.770 4.280 ;
        RECT 1001.610 4.000 1006.290 4.280 ;
        RECT 1007.130 4.000 1010.890 4.280 ;
        RECT 1011.730 4.000 1015.490 4.280 ;
        RECT 1016.330 4.000 1021.010 4.280 ;
        RECT 1021.850 4.000 1025.610 4.280 ;
        RECT 1026.450 4.000 1031.130 4.280 ;
        RECT 1031.970 4.000 1035.730 4.280 ;
        RECT 1036.570 4.000 1040.330 4.280 ;
        RECT 1041.170 4.000 1045.850 4.280 ;
        RECT 1046.690 4.000 1050.450 4.280 ;
        RECT 1051.290 4.000 1055.050 4.280 ;
        RECT 1055.890 4.000 1060.570 4.280 ;
        RECT 1061.410 4.000 1065.170 4.280 ;
        RECT 1066.010 4.000 1070.690 4.280 ;
        RECT 1071.530 4.000 1075.290 4.280 ;
        RECT 1076.130 4.000 1079.890 4.280 ;
        RECT 1080.730 4.000 1085.410 4.280 ;
        RECT 1086.250 4.000 1090.010 4.280 ;
        RECT 1090.850 4.000 1093.320 4.280 ;
      LAYER met3 ;
        RECT 4.400 1099.880 1093.905 1100.745 ;
        RECT 3.990 1093.120 1094.305 1099.880 ;
        RECT 4.400 1091.720 1093.905 1093.120 ;
        RECT 3.990 1086.320 1094.305 1091.720 ;
        RECT 4.400 1084.920 1093.905 1086.320 ;
        RECT 3.990 1079.520 1094.305 1084.920 ;
        RECT 4.400 1078.120 1093.905 1079.520 ;
        RECT 3.990 1071.360 1094.305 1078.120 ;
        RECT 4.400 1069.960 1093.905 1071.360 ;
        RECT 3.990 1064.560 1094.305 1069.960 ;
        RECT 4.400 1063.160 1093.905 1064.560 ;
        RECT 3.990 1057.760 1094.305 1063.160 ;
        RECT 4.400 1056.360 1093.905 1057.760 ;
        RECT 3.990 1049.600 1094.305 1056.360 ;
        RECT 4.400 1048.200 1093.905 1049.600 ;
        RECT 3.990 1042.800 1094.305 1048.200 ;
        RECT 4.400 1041.400 1093.905 1042.800 ;
        RECT 3.990 1034.640 1094.305 1041.400 ;
        RECT 4.400 1033.240 1093.905 1034.640 ;
        RECT 3.990 1027.840 1094.305 1033.240 ;
        RECT 4.400 1026.440 1093.905 1027.840 ;
        RECT 3.990 1021.040 1094.305 1026.440 ;
        RECT 4.400 1019.640 1093.905 1021.040 ;
        RECT 3.990 1012.880 1094.305 1019.640 ;
        RECT 4.400 1011.480 1093.905 1012.880 ;
        RECT 3.990 1006.080 1094.305 1011.480 ;
        RECT 4.400 1004.680 1093.905 1006.080 ;
        RECT 3.990 999.280 1094.305 1004.680 ;
        RECT 4.400 997.880 1093.905 999.280 ;
        RECT 3.990 991.120 1094.305 997.880 ;
        RECT 4.400 989.720 1093.905 991.120 ;
        RECT 3.990 984.320 1094.305 989.720 ;
        RECT 4.400 982.920 1093.905 984.320 ;
        RECT 3.990 976.160 1094.305 982.920 ;
        RECT 4.400 974.760 1093.905 976.160 ;
        RECT 3.990 969.360 1094.305 974.760 ;
        RECT 4.400 967.960 1093.905 969.360 ;
        RECT 3.990 962.560 1094.305 967.960 ;
        RECT 4.400 961.160 1093.905 962.560 ;
        RECT 3.990 954.400 1094.305 961.160 ;
        RECT 4.400 953.000 1093.905 954.400 ;
        RECT 3.990 947.600 1094.305 953.000 ;
        RECT 4.400 946.200 1093.905 947.600 ;
        RECT 3.990 940.800 1094.305 946.200 ;
        RECT 4.400 939.400 1093.905 940.800 ;
        RECT 3.990 932.640 1094.305 939.400 ;
        RECT 4.400 931.240 1093.905 932.640 ;
        RECT 3.990 925.840 1094.305 931.240 ;
        RECT 4.400 924.440 1093.905 925.840 ;
        RECT 3.990 917.680 1094.305 924.440 ;
        RECT 4.400 916.280 1093.905 917.680 ;
        RECT 3.990 910.880 1094.305 916.280 ;
        RECT 4.400 909.480 1093.905 910.880 ;
        RECT 3.990 904.080 1094.305 909.480 ;
        RECT 4.400 902.680 1093.905 904.080 ;
        RECT 3.990 895.920 1094.305 902.680 ;
        RECT 4.400 894.520 1093.905 895.920 ;
        RECT 3.990 889.120 1094.305 894.520 ;
        RECT 4.400 887.720 1093.905 889.120 ;
        RECT 3.990 882.320 1094.305 887.720 ;
        RECT 4.400 880.920 1093.905 882.320 ;
        RECT 3.990 874.160 1094.305 880.920 ;
        RECT 4.400 872.760 1093.905 874.160 ;
        RECT 3.990 867.360 1094.305 872.760 ;
        RECT 4.400 865.960 1093.905 867.360 ;
        RECT 3.990 859.200 1094.305 865.960 ;
        RECT 4.400 857.800 1093.905 859.200 ;
        RECT 3.990 852.400 1094.305 857.800 ;
        RECT 4.400 851.000 1093.905 852.400 ;
        RECT 3.990 845.600 1094.305 851.000 ;
        RECT 4.400 844.200 1093.905 845.600 ;
        RECT 3.990 837.440 1094.305 844.200 ;
        RECT 4.400 836.040 1093.905 837.440 ;
        RECT 3.990 830.640 1094.305 836.040 ;
        RECT 4.400 829.240 1093.905 830.640 ;
        RECT 3.990 823.840 1094.305 829.240 ;
        RECT 4.400 822.440 1093.905 823.840 ;
        RECT 3.990 815.680 1094.305 822.440 ;
        RECT 4.400 814.280 1093.905 815.680 ;
        RECT 3.990 808.880 1094.305 814.280 ;
        RECT 4.400 807.480 1093.905 808.880 ;
        RECT 3.990 800.720 1094.305 807.480 ;
        RECT 4.400 799.320 1093.905 800.720 ;
        RECT 3.990 793.920 1094.305 799.320 ;
        RECT 4.400 792.520 1093.905 793.920 ;
        RECT 3.990 787.120 1094.305 792.520 ;
        RECT 4.400 785.720 1093.905 787.120 ;
        RECT 3.990 778.960 1094.305 785.720 ;
        RECT 4.400 777.560 1093.905 778.960 ;
        RECT 3.990 772.160 1094.305 777.560 ;
        RECT 4.400 770.760 1093.905 772.160 ;
        RECT 3.990 765.360 1094.305 770.760 ;
        RECT 4.400 763.960 1093.905 765.360 ;
        RECT 3.990 757.200 1094.305 763.960 ;
        RECT 4.400 755.800 1093.905 757.200 ;
        RECT 3.990 750.400 1094.305 755.800 ;
        RECT 4.400 749.000 1093.905 750.400 ;
        RECT 3.990 742.240 1094.305 749.000 ;
        RECT 4.400 740.840 1093.905 742.240 ;
        RECT 3.990 735.440 1094.305 740.840 ;
        RECT 4.400 734.040 1093.905 735.440 ;
        RECT 3.990 728.640 1094.305 734.040 ;
        RECT 4.400 727.240 1093.905 728.640 ;
        RECT 3.990 720.480 1094.305 727.240 ;
        RECT 4.400 719.080 1093.905 720.480 ;
        RECT 3.990 713.680 1094.305 719.080 ;
        RECT 4.400 712.280 1093.905 713.680 ;
        RECT 3.990 706.880 1094.305 712.280 ;
        RECT 4.400 705.480 1093.905 706.880 ;
        RECT 3.990 698.720 1094.305 705.480 ;
        RECT 4.400 697.320 1093.905 698.720 ;
        RECT 3.990 691.920 1094.305 697.320 ;
        RECT 4.400 690.520 1093.905 691.920 ;
        RECT 3.990 683.760 1094.305 690.520 ;
        RECT 4.400 682.360 1093.905 683.760 ;
        RECT 3.990 676.960 1094.305 682.360 ;
        RECT 4.400 675.560 1093.905 676.960 ;
        RECT 3.990 670.160 1094.305 675.560 ;
        RECT 4.400 668.760 1093.905 670.160 ;
        RECT 3.990 662.000 1094.305 668.760 ;
        RECT 4.400 660.600 1093.905 662.000 ;
        RECT 3.990 655.200 1094.305 660.600 ;
        RECT 4.400 653.800 1093.905 655.200 ;
        RECT 3.990 648.400 1094.305 653.800 ;
        RECT 4.400 647.000 1093.905 648.400 ;
        RECT 3.990 640.240 1094.305 647.000 ;
        RECT 4.400 638.840 1093.905 640.240 ;
        RECT 3.990 633.440 1094.305 638.840 ;
        RECT 4.400 632.040 1093.905 633.440 ;
        RECT 3.990 625.280 1094.305 632.040 ;
        RECT 4.400 623.880 1093.905 625.280 ;
        RECT 3.990 618.480 1094.305 623.880 ;
        RECT 4.400 617.080 1093.905 618.480 ;
        RECT 3.990 611.680 1094.305 617.080 ;
        RECT 4.400 610.280 1093.905 611.680 ;
        RECT 3.990 603.520 1094.305 610.280 ;
        RECT 4.400 602.120 1093.905 603.520 ;
        RECT 3.990 596.720 1094.305 602.120 ;
        RECT 4.400 595.320 1093.905 596.720 ;
        RECT 3.990 589.920 1094.305 595.320 ;
        RECT 4.400 588.520 1093.905 589.920 ;
        RECT 3.990 581.760 1094.305 588.520 ;
        RECT 4.400 580.360 1093.905 581.760 ;
        RECT 3.990 574.960 1094.305 580.360 ;
        RECT 4.400 573.560 1093.905 574.960 ;
        RECT 3.990 566.800 1094.305 573.560 ;
        RECT 4.400 565.400 1093.905 566.800 ;
        RECT 3.990 560.000 1094.305 565.400 ;
        RECT 4.400 558.600 1093.905 560.000 ;
        RECT 3.990 553.200 1094.305 558.600 ;
        RECT 4.400 551.800 1093.905 553.200 ;
        RECT 3.990 545.040 1094.305 551.800 ;
        RECT 4.400 543.640 1093.905 545.040 ;
        RECT 3.990 538.240 1094.305 543.640 ;
        RECT 4.400 536.840 1093.905 538.240 ;
        RECT 3.990 531.440 1094.305 536.840 ;
        RECT 4.400 530.040 1093.905 531.440 ;
        RECT 3.990 523.280 1094.305 530.040 ;
        RECT 4.400 521.880 1093.905 523.280 ;
        RECT 3.990 516.480 1094.305 521.880 ;
        RECT 4.400 515.080 1093.905 516.480 ;
        RECT 3.990 508.320 1094.305 515.080 ;
        RECT 4.400 506.920 1093.905 508.320 ;
        RECT 3.990 501.520 1094.305 506.920 ;
        RECT 4.400 500.120 1093.905 501.520 ;
        RECT 3.990 494.720 1094.305 500.120 ;
        RECT 4.400 493.320 1093.905 494.720 ;
        RECT 3.990 486.560 1094.305 493.320 ;
        RECT 4.400 485.160 1093.905 486.560 ;
        RECT 3.990 479.760 1094.305 485.160 ;
        RECT 4.400 478.360 1093.905 479.760 ;
        RECT 3.990 472.960 1094.305 478.360 ;
        RECT 4.400 471.560 1093.905 472.960 ;
        RECT 3.990 464.800 1094.305 471.560 ;
        RECT 4.400 463.400 1093.905 464.800 ;
        RECT 3.990 458.000 1094.305 463.400 ;
        RECT 4.400 456.600 1093.905 458.000 ;
        RECT 3.990 449.840 1094.305 456.600 ;
        RECT 4.400 448.440 1093.905 449.840 ;
        RECT 3.990 443.040 1094.305 448.440 ;
        RECT 4.400 441.640 1093.905 443.040 ;
        RECT 3.990 436.240 1094.305 441.640 ;
        RECT 4.400 434.840 1093.905 436.240 ;
        RECT 3.990 428.080 1094.305 434.840 ;
        RECT 4.400 426.680 1093.905 428.080 ;
        RECT 3.990 421.280 1094.305 426.680 ;
        RECT 4.400 419.880 1093.905 421.280 ;
        RECT 3.990 414.480 1094.305 419.880 ;
        RECT 4.400 413.080 1093.905 414.480 ;
        RECT 3.990 406.320 1094.305 413.080 ;
        RECT 4.400 404.920 1093.905 406.320 ;
        RECT 3.990 399.520 1094.305 404.920 ;
        RECT 4.400 398.120 1093.905 399.520 ;
        RECT 3.990 391.360 1094.305 398.120 ;
        RECT 4.400 389.960 1093.905 391.360 ;
        RECT 3.990 384.560 1094.305 389.960 ;
        RECT 4.400 383.160 1093.905 384.560 ;
        RECT 3.990 377.760 1094.305 383.160 ;
        RECT 4.400 376.360 1093.905 377.760 ;
        RECT 3.990 369.600 1094.305 376.360 ;
        RECT 4.400 368.200 1093.905 369.600 ;
        RECT 3.990 362.800 1094.305 368.200 ;
        RECT 4.400 361.400 1093.905 362.800 ;
        RECT 3.990 356.000 1094.305 361.400 ;
        RECT 4.400 354.600 1093.905 356.000 ;
        RECT 3.990 347.840 1094.305 354.600 ;
        RECT 4.400 346.440 1093.905 347.840 ;
        RECT 3.990 341.040 1094.305 346.440 ;
        RECT 4.400 339.640 1093.905 341.040 ;
        RECT 3.990 332.880 1094.305 339.640 ;
        RECT 4.400 331.480 1093.905 332.880 ;
        RECT 3.990 326.080 1094.305 331.480 ;
        RECT 4.400 324.680 1093.905 326.080 ;
        RECT 3.990 319.280 1094.305 324.680 ;
        RECT 4.400 317.880 1093.905 319.280 ;
        RECT 3.990 311.120 1094.305 317.880 ;
        RECT 4.400 309.720 1093.905 311.120 ;
        RECT 3.990 304.320 1094.305 309.720 ;
        RECT 4.400 302.920 1093.905 304.320 ;
        RECT 3.990 297.520 1094.305 302.920 ;
        RECT 4.400 296.120 1093.905 297.520 ;
        RECT 3.990 289.360 1094.305 296.120 ;
        RECT 4.400 287.960 1093.905 289.360 ;
        RECT 3.990 282.560 1094.305 287.960 ;
        RECT 4.400 281.160 1093.905 282.560 ;
        RECT 3.990 274.400 1094.305 281.160 ;
        RECT 4.400 273.000 1093.905 274.400 ;
        RECT 3.990 267.600 1094.305 273.000 ;
        RECT 4.400 266.200 1093.905 267.600 ;
        RECT 3.990 260.800 1094.305 266.200 ;
        RECT 4.400 259.400 1093.905 260.800 ;
        RECT 3.990 252.640 1094.305 259.400 ;
        RECT 4.400 251.240 1093.905 252.640 ;
        RECT 3.990 245.840 1094.305 251.240 ;
        RECT 4.400 244.440 1093.905 245.840 ;
        RECT 3.990 239.040 1094.305 244.440 ;
        RECT 4.400 237.640 1093.905 239.040 ;
        RECT 3.990 230.880 1094.305 237.640 ;
        RECT 4.400 229.480 1093.905 230.880 ;
        RECT 3.990 224.080 1094.305 229.480 ;
        RECT 4.400 222.680 1093.905 224.080 ;
        RECT 3.990 215.920 1094.305 222.680 ;
        RECT 4.400 214.520 1093.905 215.920 ;
        RECT 3.990 209.120 1094.305 214.520 ;
        RECT 4.400 207.720 1093.905 209.120 ;
        RECT 3.990 202.320 1094.305 207.720 ;
        RECT 4.400 200.920 1093.905 202.320 ;
        RECT 3.990 194.160 1094.305 200.920 ;
        RECT 4.400 192.760 1093.905 194.160 ;
        RECT 3.990 187.360 1094.305 192.760 ;
        RECT 4.400 185.960 1093.905 187.360 ;
        RECT 3.990 180.560 1094.305 185.960 ;
        RECT 4.400 179.200 1094.305 180.560 ;
        RECT 4.400 179.160 1093.905 179.200 ;
        RECT 3.990 177.800 1093.905 179.160 ;
        RECT 3.990 172.400 1094.305 177.800 ;
        RECT 4.400 171.000 1093.905 172.400 ;
        RECT 3.990 165.600 1094.305 171.000 ;
        RECT 4.400 164.200 1093.905 165.600 ;
        RECT 3.990 157.440 1094.305 164.200 ;
        RECT 4.400 156.040 1093.905 157.440 ;
        RECT 3.990 150.640 1094.305 156.040 ;
        RECT 4.400 149.240 1093.905 150.640 ;
        RECT 3.990 143.840 1094.305 149.240 ;
        RECT 4.400 142.440 1093.905 143.840 ;
        RECT 3.990 135.680 1094.305 142.440 ;
        RECT 4.400 134.280 1093.905 135.680 ;
        RECT 3.990 128.880 1094.305 134.280 ;
        RECT 4.400 127.480 1093.905 128.880 ;
        RECT 3.990 122.080 1094.305 127.480 ;
        RECT 4.400 120.720 1094.305 122.080 ;
        RECT 4.400 120.680 1093.905 120.720 ;
        RECT 3.990 119.320 1093.905 120.680 ;
        RECT 3.990 113.920 1094.305 119.320 ;
        RECT 4.400 112.520 1093.905 113.920 ;
        RECT 3.990 107.120 1094.305 112.520 ;
        RECT 4.400 105.720 1093.905 107.120 ;
        RECT 3.990 98.960 1094.305 105.720 ;
        RECT 4.400 97.560 1093.905 98.960 ;
        RECT 3.990 92.160 1094.305 97.560 ;
        RECT 4.400 90.760 1093.905 92.160 ;
        RECT 3.990 85.360 1094.305 90.760 ;
        RECT 4.400 83.960 1093.905 85.360 ;
        RECT 3.990 77.200 1094.305 83.960 ;
        RECT 4.400 75.800 1093.905 77.200 ;
        RECT 3.990 70.400 1094.305 75.800 ;
        RECT 4.400 69.000 1093.905 70.400 ;
        RECT 3.990 63.600 1094.305 69.000 ;
        RECT 4.400 62.240 1094.305 63.600 ;
        RECT 4.400 62.200 1093.905 62.240 ;
        RECT 3.990 60.840 1093.905 62.200 ;
        RECT 3.990 55.440 1094.305 60.840 ;
        RECT 4.400 54.040 1093.905 55.440 ;
        RECT 3.990 48.640 1094.305 54.040 ;
        RECT 4.400 47.240 1093.905 48.640 ;
        RECT 3.990 40.480 1094.305 47.240 ;
        RECT 4.400 39.080 1093.905 40.480 ;
        RECT 3.990 33.680 1094.305 39.080 ;
        RECT 4.400 32.280 1093.905 33.680 ;
        RECT 3.990 26.880 1094.305 32.280 ;
        RECT 4.400 25.480 1093.905 26.880 ;
        RECT 3.990 18.720 1094.305 25.480 ;
        RECT 4.400 17.320 1093.905 18.720 ;
        RECT 3.990 11.920 1094.305 17.320 ;
        RECT 4.400 10.520 1093.905 11.920 ;
        RECT 3.990 4.255 1094.305 10.520 ;
      LAYER met4 ;
        RECT 15.015 10.640 1082.545 1096.400 ;
      LAYER met5 ;
        RECT 5.520 179.670 1092.500 1023.760 ;
  END
END tinyriscv
END LIBRARY

