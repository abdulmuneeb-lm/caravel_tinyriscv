magic
tech sky130A
magscale 1 2
timestamp 1609751852
<< locali >>
rect 8125 685899 8159 695453
rect 299857 666587 299891 684437
rect 364349 666587 364383 676141
rect 429577 666587 429611 684437
rect 494069 666587 494103 676141
rect 542737 666587 542771 684437
rect 299673 601715 299707 608549
rect 429393 601715 429427 608549
rect 542553 601715 542587 608549
rect 299857 589339 299891 598893
rect 429577 589339 429611 598893
rect 542737 589339 542771 598893
rect 8033 579751 8067 589237
rect 364533 550647 364567 553401
rect 429301 550647 429335 560201
rect 494253 550647 494287 553401
rect 542461 550647 542495 560201
rect 8033 540991 8067 550545
rect 299673 485775 299707 492609
rect 429393 485775 429427 492609
rect 542553 485775 542587 492609
rect 299673 466395 299707 473297
rect 429393 466395 429427 473297
rect 542553 466395 542587 473297
rect 299489 440283 299523 449837
rect 299489 423691 299523 436781
rect 8033 390575 8067 398905
rect 429301 398803 429335 405637
rect 542461 398803 542495 405637
rect 299581 389079 299615 391901
rect 364533 357527 364567 360213
rect 494253 357527 494287 360213
rect 8033 347803 8067 357357
rect 299857 356167 299891 357493
rect 8033 336855 8067 340969
rect 299857 336787 299891 354637
rect 429577 353379 429611 357493
rect 542737 353379 542771 357493
rect 364349 338147 364383 347701
rect 429669 340799 429703 353209
rect 494069 338147 494103 347701
rect 542829 340799 542863 353209
rect 7941 327131 7975 336617
rect 299673 289867 299707 299421
rect 8125 280211 8159 289765
rect 429485 280211 429519 289765
rect 542461 280211 542495 289765
rect 160109 266407 160143 266509
rect 9689 264435 9723 264537
rect 4997 261443 5031 264401
rect 19257 264367 19291 264537
rect 29009 264435 29043 264537
rect 38577 264367 38611 264537
rect 22051 264333 22109 264367
rect 41463 264333 41521 264367
rect 48329 264163 48363 264333
rect 67649 264231 67683 264333
rect 72433 264231 72467 264333
rect 81449 263823 81483 264265
rect 85589 263755 85623 264265
rect 87429 263687 87463 264265
rect 99331 264265 99389 264299
rect 89729 264163 89763 264265
rect 106289 264095 106323 264333
rect 108681 263687 108715 264265
rect 115857 264095 115891 264197
rect 133521 263891 133555 264265
rect 134441 263755 134475 264265
rect 147689 263619 147723 264265
rect 173817 263007 173851 264265
rect 202705 263823 202739 264265
rect 224417 262939 224451 264265
rect 229753 264231 229787 264333
rect 252201 263075 252235 264537
rect 259193 263619 259227 264537
rect 263609 262871 263643 266305
rect 271797 263143 271831 266237
rect 277961 264299 277995 264605
rect 278053 264435 278087 264537
rect 278697 264095 278731 264265
rect 429393 263551 429427 270453
rect 429577 253963 429611 260797
rect 429301 222207 429335 231761
rect 8033 215203 8067 222105
rect 7941 193171 7975 201433
rect 280813 200175 280847 209729
rect 280997 190859 281031 200005
rect 299673 193307 299707 202793
rect 429485 193307 429519 202793
rect 429485 173995 429519 183481
rect 429393 157335 429427 164169
rect 429393 137955 429427 144857
rect 280905 125715 280939 135201
rect 7941 115991 7975 125545
rect 280905 118643 280939 125545
rect 429301 115991 429335 125545
rect 280905 106335 280939 115889
rect 8033 99331 8067 106233
rect 280905 96679 280939 106165
rect 299673 99331 299707 101405
rect 542645 99331 542679 101405
rect 280997 89675 281031 96509
rect 280905 77299 280939 86921
rect 299673 77299 299707 86921
rect 62221 67643 62255 77197
rect 280997 67711 281031 77197
rect 280905 60639 280939 67541
rect 299673 60979 299707 67541
rect 280905 48331 280939 52717
rect 135085 38675 135119 42109
rect 137017 41327 137051 42177
rect 135085 29019 135119 38505
rect 137017 29019 137051 38573
rect 149069 37315 149103 43741
rect 146585 29019 146619 33745
rect 99205 9707 99239 27557
rect 135177 9707 135211 19193
rect 149069 18003 149103 27557
rect 150725 11679 150759 27557
rect 409797 3927 409831 4029
rect 89729 3383 89763 3485
rect 94513 3111 94547 3417
rect 101413 3247 101447 3485
rect 104173 3111 104207 3485
rect 108991 3281 109049 3315
rect 128369 3247 128403 3417
rect 425069 3383 425103 3485
rect 106289 2907 106323 3213
rect 263609 3179 263643 3349
rect 113741 2907 113775 3009
rect 152749 595 152783 2805
<< viali >>
rect 8125 695453 8159 695487
rect 8125 685865 8159 685899
rect 299857 684437 299891 684471
rect 429577 684437 429611 684471
rect 299857 666553 299891 666587
rect 364349 676141 364383 676175
rect 364349 666553 364383 666587
rect 542737 684437 542771 684471
rect 429577 666553 429611 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 542737 666553 542771 666587
rect 299673 608549 299707 608583
rect 299673 601681 299707 601715
rect 429393 608549 429427 608583
rect 429393 601681 429427 601715
rect 542553 608549 542587 608583
rect 542553 601681 542587 601715
rect 299857 598893 299891 598927
rect 299857 589305 299891 589339
rect 429577 598893 429611 598927
rect 429577 589305 429611 589339
rect 542737 598893 542771 598927
rect 542737 589305 542771 589339
rect 8033 589237 8067 589271
rect 8033 579717 8067 579751
rect 429301 560201 429335 560235
rect 364533 553401 364567 553435
rect 364533 550613 364567 550647
rect 542461 560201 542495 560235
rect 429301 550613 429335 550647
rect 494253 553401 494287 553435
rect 494253 550613 494287 550647
rect 542461 550613 542495 550647
rect 8033 550545 8067 550579
rect 8033 540957 8067 540991
rect 299673 492609 299707 492643
rect 299673 485741 299707 485775
rect 429393 492609 429427 492643
rect 429393 485741 429427 485775
rect 542553 492609 542587 492643
rect 542553 485741 542587 485775
rect 299673 473297 299707 473331
rect 299673 466361 299707 466395
rect 429393 473297 429427 473331
rect 429393 466361 429427 466395
rect 542553 473297 542587 473331
rect 542553 466361 542587 466395
rect 299489 449837 299523 449871
rect 299489 440249 299523 440283
rect 299489 436781 299523 436815
rect 299489 423657 299523 423691
rect 429301 405637 429335 405671
rect 8033 398905 8067 398939
rect 429301 398769 429335 398803
rect 542461 405637 542495 405671
rect 542461 398769 542495 398803
rect 8033 390541 8067 390575
rect 299581 391901 299615 391935
rect 299581 389045 299615 389079
rect 364533 360213 364567 360247
rect 494253 360213 494287 360247
rect 299857 357493 299891 357527
rect 364533 357493 364567 357527
rect 429577 357493 429611 357527
rect 494253 357493 494287 357527
rect 542737 357493 542771 357527
rect 8033 357357 8067 357391
rect 299857 356133 299891 356167
rect 8033 347769 8067 347803
rect 299857 354637 299891 354671
rect 8033 340969 8067 341003
rect 8033 336821 8067 336855
rect 429577 353345 429611 353379
rect 542737 353345 542771 353379
rect 429669 353209 429703 353243
rect 364349 347701 364383 347735
rect 542829 353209 542863 353243
rect 429669 340765 429703 340799
rect 494069 347701 494103 347735
rect 364349 338113 364383 338147
rect 542829 340765 542863 340799
rect 494069 338113 494103 338147
rect 299857 336753 299891 336787
rect 7941 336617 7975 336651
rect 7941 327097 7975 327131
rect 299673 299421 299707 299455
rect 299673 289833 299707 289867
rect 8125 289765 8159 289799
rect 8125 280177 8159 280211
rect 429485 289765 429519 289799
rect 429485 280177 429519 280211
rect 542461 289765 542495 289799
rect 542461 280177 542495 280211
rect 429393 270453 429427 270487
rect 160109 266509 160143 266543
rect 160109 266373 160143 266407
rect 263609 266305 263643 266339
rect 9689 264537 9723 264571
rect 4997 264401 5031 264435
rect 9689 264401 9723 264435
rect 19257 264537 19291 264571
rect 29009 264537 29043 264571
rect 29009 264401 29043 264435
rect 38577 264537 38611 264571
rect 252201 264537 252235 264571
rect 19257 264333 19291 264367
rect 22017 264333 22051 264367
rect 22109 264333 22143 264367
rect 38577 264333 38611 264367
rect 41429 264333 41463 264367
rect 41521 264333 41555 264367
rect 48329 264333 48363 264367
rect 67649 264333 67683 264367
rect 67649 264197 67683 264231
rect 72433 264333 72467 264367
rect 106289 264333 106323 264367
rect 72433 264197 72467 264231
rect 81449 264265 81483 264299
rect 48329 264129 48363 264163
rect 81449 263789 81483 263823
rect 85589 264265 85623 264299
rect 85589 263721 85623 263755
rect 87429 264265 87463 264299
rect 89729 264265 89763 264299
rect 99297 264265 99331 264299
rect 99389 264265 99423 264299
rect 89729 264129 89763 264163
rect 229753 264333 229787 264367
rect 106289 264061 106323 264095
rect 108681 264265 108715 264299
rect 87429 263653 87463 263687
rect 133521 264265 133555 264299
rect 115857 264197 115891 264231
rect 115857 264061 115891 264095
rect 133521 263857 133555 263891
rect 134441 264265 134475 264299
rect 134441 263721 134475 263755
rect 147689 264265 147723 264299
rect 108681 263653 108715 263687
rect 147689 263585 147723 263619
rect 173817 264265 173851 264299
rect 202705 264265 202739 264299
rect 202705 263789 202739 263823
rect 224417 264265 224451 264299
rect 173817 262973 173851 263007
rect 229753 264197 229787 264231
rect 259193 264537 259227 264571
rect 259193 263585 259227 263619
rect 252201 263041 252235 263075
rect 224417 262905 224451 262939
rect 271797 266237 271831 266271
rect 277961 264605 277995 264639
rect 278053 264537 278087 264571
rect 278053 264401 278087 264435
rect 277961 264265 277995 264299
rect 278697 264265 278731 264299
rect 278697 264061 278731 264095
rect 429393 263517 429427 263551
rect 271797 263109 271831 263143
rect 263609 262837 263643 262871
rect 4997 261409 5031 261443
rect 429577 260797 429611 260831
rect 429577 253929 429611 253963
rect 429301 231761 429335 231795
rect 429301 222173 429335 222207
rect 8033 222105 8067 222139
rect 8033 215169 8067 215203
rect 280813 209729 280847 209763
rect 7941 201433 7975 201467
rect 280813 200141 280847 200175
rect 299673 202793 299707 202827
rect 7941 193137 7975 193171
rect 280997 200005 281031 200039
rect 299673 193273 299707 193307
rect 429485 202793 429519 202827
rect 429485 193273 429519 193307
rect 280997 190825 281031 190859
rect 429485 183481 429519 183515
rect 429485 173961 429519 173995
rect 429393 164169 429427 164203
rect 429393 157301 429427 157335
rect 429393 144857 429427 144891
rect 429393 137921 429427 137955
rect 280905 135201 280939 135235
rect 280905 125681 280939 125715
rect 7941 125545 7975 125579
rect 280905 125545 280939 125579
rect 280905 118609 280939 118643
rect 429301 125545 429335 125579
rect 7941 115957 7975 115991
rect 429301 115957 429335 115991
rect 280905 115889 280939 115923
rect 280905 106301 280939 106335
rect 8033 106233 8067 106267
rect 8033 99297 8067 99331
rect 280905 106165 280939 106199
rect 299673 101405 299707 101439
rect 299673 99297 299707 99331
rect 542645 101405 542679 101439
rect 542645 99297 542679 99331
rect 280905 96645 280939 96679
rect 280997 96509 281031 96543
rect 280997 89641 281031 89675
rect 280905 86921 280939 86955
rect 280905 77265 280939 77299
rect 299673 86921 299707 86955
rect 299673 77265 299707 77299
rect 62221 77197 62255 77231
rect 280997 77197 281031 77231
rect 280997 67677 281031 67711
rect 62221 67609 62255 67643
rect 280905 67541 280939 67575
rect 299673 67541 299707 67575
rect 299673 60945 299707 60979
rect 280905 60605 280939 60639
rect 280905 52717 280939 52751
rect 280905 48297 280939 48331
rect 149069 43741 149103 43775
rect 137017 42177 137051 42211
rect 135085 42109 135119 42143
rect 137017 41293 137051 41327
rect 135085 38641 135119 38675
rect 137017 38573 137051 38607
rect 135085 38505 135119 38539
rect 135085 28985 135119 29019
rect 149069 37281 149103 37315
rect 137017 28985 137051 29019
rect 146585 33745 146619 33779
rect 146585 28985 146619 29019
rect 99205 27557 99239 27591
rect 149069 27557 149103 27591
rect 99205 9673 99239 9707
rect 135177 19193 135211 19227
rect 149069 17969 149103 18003
rect 150725 27557 150759 27591
rect 150725 11645 150759 11679
rect 135177 9673 135211 9707
rect 409797 4029 409831 4063
rect 409797 3893 409831 3927
rect 89729 3485 89763 3519
rect 101413 3485 101447 3519
rect 89729 3349 89763 3383
rect 94513 3417 94547 3451
rect 101413 3213 101447 3247
rect 104173 3485 104207 3519
rect 94513 3077 94547 3111
rect 425069 3485 425103 3519
rect 128369 3417 128403 3451
rect 108957 3281 108991 3315
rect 109049 3281 109083 3315
rect 104173 3077 104207 3111
rect 106289 3213 106323 3247
rect 128369 3213 128403 3247
rect 263609 3349 263643 3383
rect 425069 3349 425103 3383
rect 263609 3145 263643 3179
rect 106289 2873 106323 2907
rect 113741 3009 113775 3043
rect 113741 2873 113775 2907
rect 152749 2805 152783 2839
rect 152749 561 152783 595
<< metal1 >>
rect 111702 700680 111708 700732
rect 111760 700720 111766 700732
rect 154114 700720 154120 700732
rect 111760 700692 154120 700720
rect 111760 700680 111766 700692
rect 154114 700680 154120 700692
rect 154172 700680 154178 700732
rect 105446 700612 105452 700664
rect 105504 700652 105510 700664
rect 169754 700652 169760 700664
rect 105504 700624 169760 700652
rect 105504 700612 105510 700624
rect 169754 700612 169760 700624
rect 169812 700612 169818 700664
rect 235166 700612 235172 700664
rect 235224 700652 235230 700664
rect 235902 700652 235908 700664
rect 235224 700624 235908 700652
rect 235224 700612 235230 700624
rect 235902 700612 235908 700624
rect 235960 700612 235966 700664
rect 137830 700544 137836 700596
rect 137888 700584 137894 700596
rect 283006 700584 283012 700596
rect 137888 700556 283012 700584
rect 137888 700544 137894 700556
rect 283006 700544 283012 700556
rect 283064 700544 283070 700596
rect 72970 700476 72976 700528
rect 73028 700516 73034 700528
rect 269114 700516 269120 700528
rect 73028 700488 269120 700516
rect 73028 700476 73034 700488
rect 269114 700476 269120 700488
rect 269172 700476 269178 700528
rect 287698 700476 287704 700528
rect 287756 700516 287762 700528
rect 332502 700516 332508 700528
rect 287756 700488 332508 700516
rect 287756 700476 287762 700488
rect 332502 700476 332508 700488
rect 332560 700476 332566 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 143442 700408 143448 700460
rect 143500 700448 143506 700460
rect 348786 700448 348792 700460
rect 143500 700420 348792 700448
rect 143500 700408 143506 700420
rect 348786 700408 348792 700420
rect 348844 700408 348850 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 253934 700380 253940 700392
rect 24360 700352 253940 700380
rect 24360 700340 24366 700352
rect 253934 700340 253940 700352
rect 253992 700340 253998 700392
rect 290458 700340 290464 700392
rect 290516 700380 290522 700392
rect 413646 700380 413652 700392
rect 290516 700352 413652 700380
rect 290516 700340 290522 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 104802 700272 104808 700324
rect 104860 700312 104866 700324
rect 397454 700312 397460 700324
rect 104860 700284 397460 700312
rect 104860 700272 104866 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 399478 700272 399484 700324
rect 399536 700312 399542 700324
rect 478506 700312 478512 700324
rect 399536 700284 478512 700312
rect 399536 700272 399542 700284
rect 478506 700272 478512 700284
rect 478564 700272 478570 700324
rect 533338 700272 533344 700324
rect 533396 700312 533402 700324
rect 559650 700312 559656 700324
rect 533396 700284 559656 700312
rect 533396 700272 533402 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 542722 698232 542728 698284
rect 542780 698272 542786 698284
rect 543550 698272 543556 698284
rect 542780 698244 543556 698272
rect 542780 698232 542786 698244
rect 543550 698232 543556 698244
rect 543608 698232 543614 698284
rect 319438 696940 319444 696992
rect 319496 696980 319502 696992
rect 580166 696980 580172 696992
rect 319496 696952 580172 696980
rect 319496 696940 319502 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 282914 692792 282920 692844
rect 282972 692832 282978 692844
rect 283834 692832 283840 692844
rect 282972 692804 283840 692832
rect 282972 692792 282978 692804
rect 283834 692792 283840 692804
rect 283892 692792 283898 692844
rect 542722 688644 542728 688696
rect 542780 688644 542786 688696
rect 299658 688576 299664 688628
rect 299716 688616 299722 688628
rect 300118 688616 300124 688628
rect 299716 688588 300124 688616
rect 299716 688576 299722 688588
rect 300118 688576 300124 688588
rect 300176 688576 300182 688628
rect 429378 688576 429384 688628
rect 429436 688616 429442 688628
rect 429838 688616 429844 688628
rect 429436 688588 429844 688616
rect 429436 688576 429442 688588
rect 429838 688576 429844 688588
rect 429896 688576 429902 688628
rect 542538 688576 542544 688628
rect 542596 688616 542602 688628
rect 542740 688616 542768 688644
rect 542596 688588 542768 688616
rect 542596 688576 542602 688588
rect 299492 685936 301268 685964
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 295978 685856 295984 685908
rect 296036 685896 296042 685908
rect 299492 685896 299520 685936
rect 296036 685868 299520 685896
rect 301240 685896 301268 685936
rect 429212 685936 429976 685964
rect 429212 685896 429240 685936
rect 301240 685868 429240 685896
rect 429948 685896 429976 685936
rect 540992 685936 542860 685964
rect 540992 685896 541020 685936
rect 429948 685868 541020 685896
rect 542832 685896 542860 685936
rect 580166 685896 580172 685908
rect 542832 685868 580172 685896
rect 296036 685856 296042 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 299566 684428 299572 684480
rect 299624 684468 299630 684480
rect 299845 684471 299903 684477
rect 299845 684468 299857 684471
rect 299624 684440 299857 684468
rect 299624 684428 299630 684440
rect 299845 684437 299857 684440
rect 299891 684437 299903 684471
rect 299845 684431 299903 684437
rect 429286 684428 429292 684480
rect 429344 684468 429350 684480
rect 429565 684471 429623 684477
rect 429565 684468 429577 684471
rect 429344 684440 429577 684468
rect 429344 684428 429350 684440
rect 429565 684437 429577 684440
rect 429611 684437 429623 684471
rect 429565 684431 429623 684437
rect 542446 684428 542452 684480
rect 542504 684468 542510 684480
rect 542725 684471 542783 684477
rect 542725 684468 542737 684471
rect 542504 684440 542737 684468
rect 542504 684428 542510 684440
rect 542725 684437 542737 684440
rect 542771 684437 542783 684471
rect 542725 684431 542783 684437
rect 3326 681708 3332 681760
rect 3384 681748 3390 681760
rect 4798 681748 4804 681760
rect 3384 681720 4804 681748
rect 3384 681708 3390 681720
rect 4798 681708 4804 681720
rect 4856 681708 4862 681760
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 364334 676172 364340 676184
rect 364295 676144 364340 676172
rect 364334 676132 364340 676144
rect 364392 676132 364398 676184
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 60642 673480 60648 673532
rect 60700 673520 60706 673532
rect 580166 673520 580172 673532
rect 60700 673492 580172 673520
rect 60700 673480 60706 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 51718 667944 51724 667956
rect 3476 667916 51724 667944
rect 3476 667904 3482 667916
rect 51718 667904 51724 667916
rect 51776 667904 51782 667956
rect 299845 666587 299903 666593
rect 299845 666553 299857 666587
rect 299891 666584 299903 666587
rect 299934 666584 299940 666596
rect 299891 666556 299940 666584
rect 299891 666553 299903 666556
rect 299845 666547 299903 666553
rect 299934 666544 299940 666556
rect 299992 666544 299998 666596
rect 364337 666587 364395 666593
rect 364337 666553 364349 666587
rect 364383 666584 364395 666587
rect 364426 666584 364432 666596
rect 364383 666556 364432 666584
rect 364383 666553 364395 666556
rect 364337 666547 364395 666553
rect 364426 666544 364432 666556
rect 364484 666544 364490 666596
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 542725 666587 542783 666593
rect 542725 666553 542737 666587
rect 542771 666584 542783 666587
rect 542814 666584 542820 666596
rect 542771 666556 542820 666584
rect 542771 666553 542783 666556
rect 542725 666547 542783 666553
rect 542814 666544 542820 666556
rect 542872 666544 542878 666596
rect 8018 654100 8024 654152
rect 8076 654140 8082 654152
rect 8202 654140 8208 654152
rect 8076 654112 8208 654140
rect 8076 654100 8082 654112
rect 8202 654100 8208 654112
rect 8260 654100 8266 654152
rect 364334 654100 364340 654152
rect 364392 654140 364398 654152
rect 364518 654140 364524 654152
rect 364392 654112 364524 654140
rect 364392 654100 364398 654112
rect 364518 654100 364524 654112
rect 364576 654100 364582 654152
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 313918 650020 313924 650072
rect 313976 650060 313982 650072
rect 580166 650060 580172 650072
rect 313976 650032 580172 650060
rect 313976 650020 313982 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 299658 647232 299664 647284
rect 299716 647272 299722 647284
rect 299750 647272 299756 647284
rect 299716 647244 299756 647272
rect 299716 647232 299722 647244
rect 299750 647232 299756 647244
rect 299808 647232 299814 647284
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 542538 647232 542544 647284
rect 542596 647272 542602 647284
rect 542630 647272 542636 647284
rect 542596 647244 542636 647272
rect 542596 647232 542602 647244
rect 542630 647232 542636 647244
rect 542688 647232 542694 647284
rect 299658 640364 299664 640416
rect 299716 640404 299722 640416
rect 299750 640404 299756 640416
rect 299716 640376 299756 640404
rect 299716 640364 299722 640376
rect 299750 640364 299756 640376
rect 299808 640364 299814 640416
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 542538 640364 542544 640416
rect 542596 640404 542602 640416
rect 542630 640404 542636 640416
rect 542596 640376 542636 640404
rect 542596 640364 542602 640376
rect 542630 640364 542636 640376
rect 542688 640364 542694 640416
rect 293218 638936 293224 638988
rect 293276 638976 293282 638988
rect 580166 638976 580172 638988
rect 293276 638948 580172 638976
rect 293276 638936 293282 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 8018 634788 8024 634840
rect 8076 634828 8082 634840
rect 8202 634828 8208 634840
rect 8076 634800 8208 634828
rect 8076 634788 8082 634800
rect 8202 634788 8208 634800
rect 8260 634788 8266 634840
rect 364334 634788 364340 634840
rect 364392 634828 364398 634840
rect 364518 634828 364524 634840
rect 364392 634800 364524 634828
rect 364392 634788 364398 634800
rect 364518 634788 364524 634800
rect 364576 634788 364582 634840
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 299566 630640 299572 630692
rect 299624 630680 299630 630692
rect 299750 630680 299756 630692
rect 299624 630652 299756 630680
rect 299624 630640 299630 630652
rect 299750 630640 299756 630652
rect 299808 630640 299814 630692
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 542446 630640 542452 630692
rect 542504 630680 542510 630692
rect 542630 630680 542636 630692
rect 542504 630652 542636 630680
rect 542504 630640 542510 630652
rect 542630 630640 542636 630652
rect 542688 630640 542694 630692
rect 284938 626560 284944 626612
rect 284996 626600 285002 626612
rect 580166 626600 580172 626612
rect 284996 626572 580172 626600
rect 284996 626560 285002 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 4062 623772 4068 623824
rect 4120 623812 4126 623824
rect 6178 623812 6184 623824
rect 4120 623784 6184 623812
rect 4120 623772 4126 623784
rect 6178 623772 6184 623784
rect 6236 623772 6242 623824
rect 8018 615476 8024 615528
rect 8076 615516 8082 615528
rect 8202 615516 8208 615528
rect 8076 615488 8208 615516
rect 8076 615476 8082 615488
rect 8202 615476 8208 615488
rect 8260 615476 8266 615528
rect 364334 615476 364340 615528
rect 364392 615516 364398 615528
rect 364518 615516 364524 615528
rect 364392 615488 364524 615516
rect 364392 615476 364398 615488
rect 364518 615476 364524 615488
rect 364576 615476 364582 615528
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 299566 611328 299572 611380
rect 299624 611368 299630 611380
rect 299750 611368 299756 611380
rect 299624 611340 299756 611368
rect 299624 611328 299630 611340
rect 299750 611328 299756 611340
rect 299808 611328 299814 611380
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 542446 611328 542452 611380
rect 542504 611368 542510 611380
rect 542630 611368 542636 611380
rect 542504 611340 542636 611368
rect 542504 611328 542510 611340
rect 542630 611328 542636 611340
rect 542688 611328 542694 611380
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 14550 610008 14556 610020
rect 3476 609980 14556 610008
rect 3476 609968 3482 609980
rect 14550 609968 14556 609980
rect 14608 609968 14614 610020
rect 299658 608580 299664 608592
rect 299619 608552 299664 608580
rect 299658 608540 299664 608552
rect 299716 608540 299722 608592
rect 429378 608580 429384 608592
rect 429339 608552 429384 608580
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 542538 608580 542544 608592
rect 542499 608552 542544 608580
rect 542538 608540 542544 608552
rect 542596 608540 542602 608592
rect 223482 603100 223488 603152
rect 223540 603140 223546 603152
rect 580166 603140 580172 603152
rect 223540 603112 580172 603140
rect 223540 603100 223546 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 299661 601715 299719 601721
rect 299661 601681 299673 601715
rect 299707 601712 299719 601715
rect 299842 601712 299848 601724
rect 299707 601684 299848 601712
rect 299707 601681 299719 601684
rect 299661 601675 299719 601681
rect 299842 601672 299848 601684
rect 299900 601672 299906 601724
rect 429381 601715 429439 601721
rect 429381 601681 429393 601715
rect 429427 601712 429439 601715
rect 429562 601712 429568 601724
rect 429427 601684 429568 601712
rect 429427 601681 429439 601684
rect 429381 601675 429439 601681
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 542541 601715 542599 601721
rect 542541 601681 542553 601715
rect 542587 601712 542599 601715
rect 542722 601712 542728 601724
rect 542587 601684 542728 601712
rect 542587 601681 542599 601684
rect 542541 601675 542599 601681
rect 542722 601672 542728 601684
rect 542780 601672 542786 601724
rect 299842 598924 299848 598936
rect 299803 598896 299848 598924
rect 299842 598884 299848 598896
rect 299900 598884 299906 598936
rect 429562 598924 429568 598936
rect 429523 598896 429568 598924
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 542722 598924 542728 598936
rect 542683 598896 542728 598924
rect 542722 598884 542728 598896
rect 542780 598884 542786 598936
rect 8018 596164 8024 596216
rect 8076 596204 8082 596216
rect 8202 596204 8208 596216
rect 8076 596176 8208 596204
rect 8076 596164 8082 596176
rect 8202 596164 8208 596176
rect 8260 596164 8266 596216
rect 364334 596164 364340 596216
rect 364392 596204 364398 596216
rect 364518 596204 364524 596216
rect 364392 596176 364524 596204
rect 364392 596164 364398 596176
rect 364518 596164 364524 596176
rect 364576 596164 364582 596216
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 190454 594844 190460 594856
rect 3292 594816 190460 594844
rect 3292 594804 3298 594816
rect 190454 594804 190460 594816
rect 190512 594804 190518 594856
rect 73062 592016 73068 592068
rect 73120 592056 73126 592068
rect 580166 592056 580172 592068
rect 73120 592028 580172 592056
rect 73120 592016 73126 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 299845 589339 299903 589345
rect 299845 589305 299857 589339
rect 299891 589336 299903 589339
rect 299934 589336 299940 589348
rect 299891 589308 299940 589336
rect 299891 589305 299903 589308
rect 299845 589299 299903 589305
rect 299934 589296 299940 589308
rect 299992 589296 299998 589348
rect 429565 589339 429623 589345
rect 429565 589305 429577 589339
rect 429611 589336 429623 589339
rect 429654 589336 429660 589348
rect 429611 589308 429660 589336
rect 429611 589305 429623 589308
rect 429565 589299 429623 589305
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 542725 589339 542783 589345
rect 542725 589305 542737 589339
rect 542771 589336 542783 589339
rect 542814 589336 542820 589348
rect 542771 589308 542820 589336
rect 542771 589305 542783 589308
rect 542725 589299 542783 589305
rect 542814 589296 542820 589308
rect 542872 589296 542878 589348
rect 8018 589268 8024 589280
rect 7979 589240 8024 589268
rect 8018 589228 8024 589240
rect 8076 589228 8082 589280
rect 364150 589228 364156 589280
rect 364208 589268 364214 589280
rect 364426 589268 364432 589280
rect 364208 589240 364432 589268
rect 364208 589228 364214 589240
rect 364426 589228 364432 589240
rect 364484 589228 364490 589280
rect 493870 589228 493876 589280
rect 493928 589268 493934 589280
rect 494146 589268 494152 589280
rect 493928 589240 494152 589268
rect 493928 589228 493934 589240
rect 494146 589228 494152 589240
rect 494204 589228 494210 589280
rect 299934 582468 299940 582480
rect 299860 582440 299940 582468
rect 299860 582344 299888 582440
rect 299934 582428 299940 582440
rect 299992 582428 299998 582480
rect 429654 582468 429660 582480
rect 429580 582440 429660 582468
rect 429580 582344 429608 582440
rect 429654 582428 429660 582440
rect 429712 582428 429718 582480
rect 542814 582468 542820 582480
rect 542740 582440 542820 582468
rect 542740 582344 542768 582440
rect 542814 582428 542820 582440
rect 542872 582428 542878 582480
rect 299842 582292 299848 582344
rect 299900 582292 299906 582344
rect 429562 582292 429568 582344
rect 429620 582292 429626 582344
rect 542722 582292 542728 582344
rect 542780 582292 542786 582344
rect 8018 579748 8024 579760
rect 7979 579720 8024 579748
rect 8018 579708 8024 579720
rect 8076 579708 8082 579760
rect 329098 579640 329104 579692
rect 329156 579680 329162 579692
rect 580166 579680 580172 579692
rect 329156 579652 580172 579680
rect 329156 579640 329162 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 7926 579572 7932 579624
rect 7984 579612 7990 579624
rect 8110 579612 8116 579624
rect 7984 579584 8116 579612
rect 7984 579572 7990 579584
rect 8110 579572 8116 579584
rect 8168 579572 8174 579624
rect 4062 567196 4068 567248
rect 4120 567236 4126 567248
rect 255314 567236 255320 567248
rect 4120 567208 255320 567236
rect 4120 567196 4126 567208
rect 255314 567196 255320 567208
rect 255372 567196 255378 567248
rect 429286 563116 429292 563168
rect 429344 563116 429350 563168
rect 542446 563116 542452 563168
rect 542504 563116 542510 563168
rect 429304 563032 429332 563116
rect 542464 563032 542492 563116
rect 429286 562980 429292 563032
rect 429344 562980 429350 563032
rect 542446 562980 542452 563032
rect 542504 562980 542510 563032
rect 7926 562912 7932 562964
rect 7984 562952 7990 562964
rect 8110 562952 8116 562964
rect 7984 562924 8116 562952
rect 7984 562912 7990 562924
rect 8110 562912 8116 562924
rect 8168 562912 8174 562964
rect 429286 560232 429292 560244
rect 429247 560204 429292 560232
rect 429286 560192 429292 560204
rect 429344 560192 429350 560244
rect 542446 560232 542452 560244
rect 542407 560204 542452 560232
rect 542446 560192 542452 560204
rect 542504 560192 542510 560244
rect 521654 556384 521660 556436
rect 521712 556424 521718 556436
rect 529290 556424 529296 556436
rect 521712 556396 529296 556424
rect 521712 556384 521718 556396
rect 529290 556384 529296 556396
rect 529348 556384 529354 556436
rect 415394 556316 415400 556368
rect 415452 556356 415458 556368
rect 424870 556356 424876 556368
rect 415452 556328 424876 556356
rect 415452 556316 415458 556328
rect 424870 556316 424876 556328
rect 424928 556316 424934 556368
rect 364518 553432 364524 553444
rect 364479 553404 364524 553432
rect 364518 553392 364524 553404
rect 364576 553392 364582 553444
rect 494238 553432 494244 553444
rect 494199 553404 494244 553432
rect 494238 553392 494244 553404
rect 494296 553392 494302 553444
rect 4062 552032 4068 552084
rect 4120 552072 4126 552084
rect 15838 552072 15844 552084
rect 4120 552044 15844 552072
rect 4120 552032 4126 552044
rect 15838 552032 15844 552044
rect 15896 552032 15902 552084
rect 299474 550604 299480 550656
rect 299532 550644 299538 550656
rect 299658 550644 299664 550656
rect 299532 550616 299664 550644
rect 299532 550604 299538 550616
rect 299658 550604 299664 550616
rect 299716 550604 299722 550656
rect 364518 550644 364524 550656
rect 364479 550616 364524 550644
rect 364518 550604 364524 550616
rect 364576 550604 364582 550656
rect 429289 550647 429347 550653
rect 429289 550613 429301 550647
rect 429335 550644 429347 550647
rect 429470 550644 429476 550656
rect 429335 550616 429476 550644
rect 429335 550613 429347 550616
rect 429289 550607 429347 550613
rect 429470 550604 429476 550616
rect 429528 550604 429534 550656
rect 494238 550644 494244 550656
rect 494199 550616 494244 550644
rect 494238 550604 494244 550616
rect 494296 550604 494302 550656
rect 542449 550647 542507 550653
rect 542449 550613 542461 550647
rect 542495 550644 542507 550647
rect 542630 550644 542636 550656
rect 542495 550616 542636 550644
rect 542495 550613 542507 550616
rect 542449 550607 542507 550613
rect 542630 550604 542636 550616
rect 542688 550604 542694 550656
rect 8018 550576 8024 550588
rect 7979 550548 8024 550576
rect 8018 550536 8024 550548
rect 8076 550536 8082 550588
rect 281442 545096 281448 545148
rect 281500 545136 281506 545148
rect 580166 545136 580172 545148
rect 281500 545108 580172 545136
rect 281500 545096 281506 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 364518 543804 364524 543856
rect 364576 543804 364582 543856
rect 494238 543804 494244 543856
rect 494296 543804 494302 543856
rect 364536 543776 364564 543804
rect 364610 543776 364616 543788
rect 364536 543748 364616 543776
rect 364610 543736 364616 543748
rect 364668 543736 364674 543788
rect 494256 543776 494284 543804
rect 494330 543776 494336 543788
rect 494256 543748 494336 543776
rect 494330 543736 494336 543748
rect 494388 543736 494394 543788
rect 299290 543668 299296 543720
rect 299348 543708 299354 543720
rect 299474 543708 299480 543720
rect 299348 543680 299480 543708
rect 299348 543668 299354 543680
rect 299474 543668 299480 543680
rect 299532 543668 299538 543720
rect 429286 543600 429292 543652
rect 429344 543640 429350 543652
rect 429470 543640 429476 543652
rect 429344 543612 429476 543640
rect 429344 543600 429350 543612
rect 429470 543600 429476 543612
rect 429528 543600 429534 543652
rect 542446 543600 542452 543652
rect 542504 543640 542510 543652
rect 542630 543640 542636 543652
rect 542504 543612 542636 543640
rect 542504 543600 542510 543612
rect 542630 543600 542636 543612
rect 542688 543600 542694 543652
rect 8021 540991 8079 540997
rect 8021 540957 8033 540991
rect 8067 540988 8079 540991
rect 8202 540988 8208 541000
rect 8067 540960 8208 540988
rect 8067 540957 8079 540960
rect 8021 540951 8079 540957
rect 8202 540948 8208 540960
rect 8260 540948 8266 541000
rect 3970 538432 3976 538484
rect 4028 538472 4034 538484
rect 10318 538472 10324 538484
rect 4028 538444 10324 538472
rect 4028 538432 4034 538444
rect 10318 538432 10324 538444
rect 10376 538432 10382 538484
rect 429286 534012 429292 534064
rect 429344 534052 429350 534064
rect 429470 534052 429476 534064
rect 429344 534024 429476 534052
rect 429344 534012 429350 534024
rect 429470 534012 429476 534024
rect 429528 534012 429534 534064
rect 542446 534012 542452 534064
rect 542504 534052 542510 534064
rect 542630 534052 542636 534064
rect 542504 534024 542636 534052
rect 542504 534012 542510 534024
rect 542630 534012 542636 534024
rect 542688 534012 542694 534064
rect 249702 532720 249708 532772
rect 249760 532760 249766 532772
rect 580166 532760 580172 532772
rect 249760 532732 580172 532760
rect 249760 532720 249766 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 299566 531292 299572 531344
rect 299624 531332 299630 531344
rect 299750 531332 299756 531344
rect 299624 531304 299756 531332
rect 299624 531292 299630 531304
rect 299750 531292 299756 531304
rect 299808 531292 299814 531344
rect 364426 531292 364432 531344
rect 364484 531332 364490 531344
rect 364702 531332 364708 531344
rect 364484 531304 364708 531332
rect 364484 531292 364490 531304
rect 364702 531292 364708 531304
rect 364760 531292 364766 531344
rect 494146 531292 494152 531344
rect 494204 531332 494210 531344
rect 494422 531332 494428 531344
rect 494204 531304 494428 531332
rect 494204 531292 494210 531304
rect 494422 531292 494428 531304
rect 494480 531292 494486 531344
rect 364702 524532 364708 524544
rect 364628 524504 364708 524532
rect 299750 524424 299756 524476
rect 299808 524424 299814 524476
rect 299768 524396 299796 524424
rect 364628 524408 364656 524504
rect 364702 524492 364708 524504
rect 364760 524492 364766 524544
rect 494422 524532 494428 524544
rect 494348 524504 494428 524532
rect 429470 524424 429476 524476
rect 429528 524424 429534 524476
rect 299842 524396 299848 524408
rect 299768 524368 299848 524396
rect 299842 524356 299848 524368
rect 299900 524356 299906 524408
rect 364610 524356 364616 524408
rect 364668 524356 364674 524408
rect 429488 524396 429516 524424
rect 494348 524408 494376 524504
rect 494422 524492 494428 524504
rect 494480 524492 494486 524544
rect 542630 524424 542636 524476
rect 542688 524424 542694 524476
rect 429562 524396 429568 524408
rect 429488 524368 429568 524396
rect 429562 524356 429568 524368
rect 429620 524356 429626 524408
rect 494330 524356 494336 524408
rect 494388 524356 494394 524408
rect 542648 524396 542676 524424
rect 542722 524396 542728 524408
rect 542648 524368 542728 524396
rect 542722 524356 542728 524368
rect 542780 524356 542786 524408
rect 8202 521636 8208 521688
rect 8260 521676 8266 521688
rect 8386 521676 8392 521688
rect 8260 521648 8392 521676
rect 8260 521636 8266 521648
rect 8386 521636 8392 521648
rect 8444 521636 8450 521688
rect 299658 511980 299664 512032
rect 299716 512020 299722 512032
rect 299934 512020 299940 512032
rect 299716 511992 299940 512020
rect 299716 511980 299722 511992
rect 299934 511980 299940 511992
rect 299992 511980 299998 512032
rect 364426 511980 364432 512032
rect 364484 512020 364490 512032
rect 364702 512020 364708 512032
rect 364484 511992 364708 512020
rect 364484 511980 364490 511992
rect 364702 511980 364708 511992
rect 364760 511980 364766 512032
rect 429378 511980 429384 512032
rect 429436 512020 429442 512032
rect 429654 512020 429660 512032
rect 429436 511992 429660 512020
rect 429436 511980 429442 511992
rect 429654 511980 429660 511992
rect 429712 511980 429718 512032
rect 494146 511980 494152 512032
rect 494204 512020 494210 512032
rect 494422 512020 494428 512032
rect 494204 511992 494428 512020
rect 494204 511980 494210 511992
rect 494422 511980 494428 511992
rect 494480 511980 494486 512032
rect 542538 511980 542544 512032
rect 542596 512020 542602 512032
rect 542814 512020 542820 512032
rect 542596 511992 542820 512020
rect 542596 511980 542602 511992
rect 542814 511980 542820 511992
rect 542872 511980 542878 512032
rect 3878 509260 3884 509312
rect 3936 509300 3942 509312
rect 242894 509300 242900 509312
rect 3936 509272 242900 509300
rect 3936 509260 3942 509272
rect 242894 509260 242900 509272
rect 242952 509260 242958 509312
rect 285030 509260 285036 509312
rect 285088 509300 285094 509312
rect 580166 509300 580172 509312
rect 285088 509272 580172 509300
rect 285088 509260 285094 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 8202 502324 8208 502376
rect 8260 502364 8266 502376
rect 8386 502364 8392 502376
rect 8260 502336 8392 502364
rect 8260 502324 8266 502336
rect 8386 502324 8392 502336
rect 8444 502324 8450 502376
rect 299750 502324 299756 502376
rect 299808 502364 299814 502376
rect 299934 502364 299940 502376
rect 299808 502336 299940 502364
rect 299808 502324 299814 502336
rect 299934 502324 299940 502336
rect 299992 502324 299998 502376
rect 364518 502324 364524 502376
rect 364576 502364 364582 502376
rect 364702 502364 364708 502376
rect 364576 502336 364708 502364
rect 364576 502324 364582 502336
rect 364702 502324 364708 502336
rect 364760 502324 364766 502376
rect 429470 502324 429476 502376
rect 429528 502364 429534 502376
rect 429654 502364 429660 502376
rect 429528 502336 429660 502364
rect 429528 502324 429534 502336
rect 429654 502324 429660 502336
rect 429712 502324 429718 502376
rect 494238 502324 494244 502376
rect 494296 502364 494302 502376
rect 494422 502364 494428 502376
rect 494296 502336 494428 502364
rect 494296 502324 494302 502336
rect 494422 502324 494428 502336
rect 494480 502324 494486 502376
rect 542630 502324 542636 502376
rect 542688 502364 542694 502376
rect 542814 502364 542820 502376
rect 542688 502336 542820 502364
rect 542688 502324 542694 502336
rect 542814 502324 542820 502336
rect 542872 502324 542878 502376
rect 294598 498176 294604 498228
rect 294656 498216 294662 498228
rect 580166 498216 580172 498228
rect 294656 498188 580172 498216
rect 294656 498176 294662 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 4062 495456 4068 495508
rect 4120 495496 4126 495508
rect 205634 495496 205640 495508
rect 4120 495468 205640 495496
rect 4120 495456 4126 495468
rect 205634 495456 205640 495468
rect 205692 495456 205698 495508
rect 7926 492600 7932 492652
rect 7984 492640 7990 492652
rect 8110 492640 8116 492652
rect 7984 492612 8116 492640
rect 7984 492600 7990 492612
rect 8110 492600 8116 492612
rect 8168 492600 8174 492652
rect 299658 492640 299664 492652
rect 299619 492612 299664 492640
rect 299658 492600 299664 492612
rect 299716 492600 299722 492652
rect 429378 492640 429384 492652
rect 429339 492612 429384 492640
rect 429378 492600 429384 492612
rect 429436 492600 429442 492652
rect 542538 492640 542544 492652
rect 542499 492612 542544 492640
rect 542538 492600 542544 492612
rect 542596 492600 542602 492652
rect 291838 485800 291844 485852
rect 291896 485840 291902 485852
rect 580166 485840 580172 485852
rect 291896 485812 580172 485840
rect 291896 485800 291902 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 299658 485772 299664 485784
rect 299619 485744 299664 485772
rect 299658 485732 299664 485744
rect 299716 485732 299722 485784
rect 429378 485772 429384 485784
rect 429339 485744 429384 485772
rect 429378 485732 429384 485744
rect 429436 485732 429442 485784
rect 542538 485772 542544 485784
rect 542499 485744 542544 485772
rect 542538 485732 542544 485744
rect 542596 485732 542602 485784
rect 3326 480564 3332 480616
rect 3384 480604 3390 480616
rect 11698 480604 11704 480616
rect 3384 480576 11704 480604
rect 3384 480564 3390 480576
rect 11698 480564 11704 480576
rect 11756 480564 11762 480616
rect 364334 480224 364340 480276
rect 364392 480264 364398 480276
rect 364518 480264 364524 480276
rect 364392 480236 364524 480264
rect 364392 480224 364398 480236
rect 364518 480224 364524 480236
rect 364576 480224 364582 480276
rect 494054 480224 494060 480276
rect 494112 480264 494118 480276
rect 494238 480264 494244 480276
rect 494112 480236 494244 480264
rect 494112 480224 494118 480236
rect 494238 480224 494244 480236
rect 494296 480224 494302 480276
rect 299566 476076 299572 476128
rect 299624 476116 299630 476128
rect 299750 476116 299756 476128
rect 299624 476088 299756 476116
rect 299624 476076 299630 476088
rect 299750 476076 299756 476088
rect 299808 476076 299814 476128
rect 429286 476076 429292 476128
rect 429344 476116 429350 476128
rect 429470 476116 429476 476128
rect 429344 476088 429476 476116
rect 429344 476076 429350 476088
rect 429470 476076 429476 476088
rect 429528 476076 429534 476128
rect 542446 476076 542452 476128
rect 542504 476116 542510 476128
rect 542630 476116 542636 476128
rect 542504 476088 542636 476116
rect 542504 476076 542510 476088
rect 542630 476076 542636 476088
rect 542688 476076 542694 476128
rect 8018 473288 8024 473340
rect 8076 473328 8082 473340
rect 8110 473328 8116 473340
rect 8076 473300 8116 473328
rect 8076 473288 8082 473300
rect 8110 473288 8116 473300
rect 8168 473288 8174 473340
rect 299658 473328 299664 473340
rect 299619 473300 299664 473328
rect 299658 473288 299664 473300
rect 299716 473288 299722 473340
rect 429378 473328 429384 473340
rect 429339 473300 429384 473328
rect 429378 473288 429384 473300
rect 429436 473288 429442 473340
rect 542538 473328 542544 473340
rect 542499 473300 542544 473328
rect 542538 473288 542544 473300
rect 542596 473288 542602 473340
rect 299658 466392 299664 466404
rect 299619 466364 299664 466392
rect 299658 466352 299664 466364
rect 299716 466352 299722 466404
rect 429378 466392 429384 466404
rect 429339 466364 429384 466392
rect 429378 466352 429384 466364
rect 429436 466352 429442 466404
rect 542538 466392 542544 466404
rect 542499 466364 542544 466392
rect 542538 466352 542544 466364
rect 542596 466352 542602 466404
rect 160002 462340 160008 462392
rect 160060 462380 160066 462392
rect 580166 462380 580172 462392
rect 160060 462352 580172 462380
rect 160060 462340 160066 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 235902 461592 235908 461644
rect 235960 461632 235966 461644
rect 281534 461632 281540 461644
rect 235960 461604 281540 461632
rect 235960 461592 235966 461604
rect 281534 461592 281540 461604
rect 281592 461592 281598 461644
rect 364334 460912 364340 460964
rect 364392 460952 364398 460964
rect 364518 460952 364524 460964
rect 364392 460924 364524 460952
rect 364392 460912 364398 460924
rect 364518 460912 364524 460924
rect 364576 460912 364582 460964
rect 494054 460912 494060 460964
rect 494112 460952 494118 460964
rect 494238 460952 494244 460964
rect 494112 460924 494244 460952
rect 494112 460912 494118 460924
rect 494238 460912 494244 460924
rect 494296 460912 494302 460964
rect 299382 460844 299388 460896
rect 299440 460884 299446 460896
rect 299750 460884 299756 460896
rect 299440 460856 299756 460884
rect 299440 460844 299446 460856
rect 299750 460844 299756 460856
rect 299808 460844 299814 460896
rect 299400 451336 299888 451364
rect 100662 451256 100668 451308
rect 100720 451296 100726 451308
rect 299400 451296 299428 451336
rect 100720 451268 299428 451296
rect 299860 451296 299888 451336
rect 580166 451296 580172 451308
rect 299860 451268 580172 451296
rect 100720 451256 100726 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 299474 449868 299480 449880
rect 299435 449840 299480 449868
rect 299474 449828 299480 449840
rect 299532 449828 299538 449880
rect 8018 447108 8024 447160
rect 8076 447108 8082 447160
rect 429194 447108 429200 447160
rect 429252 447108 429258 447160
rect 542354 447108 542360 447160
rect 542412 447108 542418 447160
rect 8036 447080 8064 447108
rect 8110 447080 8116 447092
rect 8036 447052 8116 447080
rect 8110 447040 8116 447052
rect 8168 447040 8174 447092
rect 429212 447080 429240 447108
rect 429286 447080 429292 447092
rect 429212 447052 429292 447080
rect 429286 447040 429292 447052
rect 429344 447040 429350 447092
rect 542372 447080 542400 447108
rect 542446 447080 542452 447092
rect 542372 447052 542452 447080
rect 542446 447040 542452 447052
rect 542504 447040 542510 447092
rect 7834 444320 7840 444372
rect 7892 444360 7898 444372
rect 8110 444360 8116 444372
rect 7892 444332 8116 444360
rect 7892 444320 7898 444332
rect 8110 444320 8116 444332
rect 8168 444320 8174 444372
rect 429010 444320 429016 444372
rect 429068 444360 429074 444372
rect 429286 444360 429292 444372
rect 429068 444332 429292 444360
rect 429068 444320 429074 444332
rect 429286 444320 429292 444332
rect 429344 444320 429350 444372
rect 542170 444320 542176 444372
rect 542228 444360 542234 444372
rect 542446 444360 542452 444372
rect 542228 444332 542452 444360
rect 542228 444320 542234 444332
rect 542446 444320 542452 444332
rect 542504 444320 542510 444372
rect 364334 441600 364340 441652
rect 364392 441640 364398 441652
rect 364518 441640 364524 441652
rect 364392 441612 364524 441640
rect 364392 441600 364398 441612
rect 364518 441600 364524 441612
rect 364576 441600 364582 441652
rect 494054 441600 494060 441652
rect 494112 441640 494118 441652
rect 494238 441640 494244 441652
rect 494112 441612 494244 441640
rect 494112 441600 494118 441612
rect 494238 441600 494244 441612
rect 494296 441600 494302 441652
rect 299477 440283 299535 440289
rect 299477 440249 299489 440283
rect 299523 440280 299535 440283
rect 299566 440280 299572 440292
rect 299523 440252 299572 440280
rect 299523 440249 299535 440252
rect 299477 440243 299535 440249
rect 299566 440240 299572 440252
rect 299624 440240 299630 440292
rect 62482 438880 62488 438932
rect 62540 438920 62546 438932
rect 580166 438920 580172 438932
rect 62540 438892 580172 438920
rect 62540 438880 62546 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 3786 437452 3792 437504
rect 3844 437492 3850 437504
rect 14458 437492 14464 437504
rect 3844 437464 14464 437492
rect 3844 437452 3850 437464
rect 14458 437452 14464 437464
rect 14516 437452 14522 437504
rect 299477 436815 299535 436821
rect 299477 436781 299489 436815
rect 299523 436812 299535 436815
rect 299566 436812 299572 436824
rect 299523 436784 299572 436812
rect 299523 436781 299535 436784
rect 299477 436775 299535 436781
rect 299566 436772 299572 436784
rect 299624 436772 299630 436824
rect 8018 427864 8024 427916
rect 8076 427864 8082 427916
rect 8036 427780 8064 427864
rect 429194 427796 429200 427848
rect 429252 427796 429258 427848
rect 542354 427796 542360 427848
rect 542412 427796 542418 427848
rect 8018 427728 8024 427780
rect 8076 427728 8082 427780
rect 429212 427768 429240 427796
rect 429286 427768 429292 427780
rect 429212 427740 429292 427768
rect 429286 427728 429292 427740
rect 429344 427728 429350 427780
rect 542372 427768 542400 427796
rect 542446 427768 542452 427780
rect 542372 427740 542452 427768
rect 542446 427728 542452 427740
rect 542504 427728 542510 427780
rect 429010 425008 429016 425060
rect 429068 425048 429074 425060
rect 429286 425048 429292 425060
rect 429068 425020 429292 425048
rect 429068 425008 429074 425020
rect 429286 425008 429292 425020
rect 429344 425008 429350 425060
rect 542170 425008 542176 425060
rect 542228 425048 542234 425060
rect 542446 425048 542452 425060
rect 542228 425020 542452 425048
rect 542228 425008 542234 425020
rect 542446 425008 542452 425020
rect 542504 425008 542510 425060
rect 4062 423648 4068 423700
rect 4120 423688 4126 423700
rect 13078 423688 13084 423700
rect 4120 423660 13084 423688
rect 4120 423648 4126 423660
rect 13078 423648 13084 423660
rect 13136 423648 13142 423700
rect 299477 423691 299535 423697
rect 299477 423657 299489 423691
rect 299523 423688 299535 423691
rect 299566 423688 299572 423700
rect 299523 423660 299572 423688
rect 299523 423657 299535 423660
rect 299477 423651 299535 423657
rect 299566 423648 299572 423660
rect 299624 423648 299630 423700
rect 364334 422288 364340 422340
rect 364392 422328 364398 422340
rect 364518 422328 364524 422340
rect 364392 422300 364524 422328
rect 364392 422288 364398 422300
rect 364518 422288 364524 422300
rect 364576 422288 364582 422340
rect 494054 422288 494060 422340
rect 494112 422328 494118 422340
rect 494238 422328 494244 422340
rect 494112 422300 494244 422328
rect 494112 422288 494118 422300
rect 494238 422288 494244 422300
rect 494296 422288 494302 422340
rect 299566 422220 299572 422272
rect 299624 422260 299630 422272
rect 299750 422260 299756 422272
rect 299624 422232 299756 422260
rect 299624 422220 299630 422232
rect 299750 422220 299756 422232
rect 299808 422220 299814 422272
rect 8018 418140 8024 418192
rect 8076 418180 8082 418192
rect 8202 418180 8208 418192
rect 8076 418152 8208 418180
rect 8076 418140 8082 418152
rect 8202 418140 8208 418152
rect 8260 418140 8266 418192
rect 315298 415420 315304 415472
rect 315356 415460 315362 415472
rect 580166 415460 580172 415472
rect 315356 415432 580172 415460
rect 315356 415420 315362 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 299474 412564 299480 412616
rect 299532 412604 299538 412616
rect 299566 412604 299572 412616
rect 299532 412576 299572 412604
rect 299532 412564 299538 412576
rect 299566 412564 299572 412576
rect 299624 412564 299630 412616
rect 429194 408484 429200 408536
rect 429252 408484 429258 408536
rect 542354 408484 542360 408536
rect 542412 408484 542418 408536
rect 429212 408388 429240 408484
rect 429286 408388 429292 408400
rect 429212 408360 429292 408388
rect 429286 408348 429292 408360
rect 429344 408348 429350 408400
rect 542372 408388 542400 408484
rect 542446 408388 542452 408400
rect 542372 408360 542452 408388
rect 542446 408348 542452 408360
rect 542504 408348 542510 408400
rect 429286 405668 429292 405680
rect 429247 405640 429292 405668
rect 429286 405628 429292 405640
rect 429344 405628 429350 405680
rect 542446 405668 542452 405680
rect 542407 405640 542452 405668
rect 542446 405628 542452 405640
rect 542504 405628 542510 405680
rect 286318 404336 286324 404388
rect 286376 404376 286382 404388
rect 580166 404376 580172 404388
rect 286376 404348 580172 404376
rect 286376 404336 286382 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 364334 402976 364340 403028
rect 364392 403016 364398 403028
rect 364518 403016 364524 403028
rect 364392 402988 364524 403016
rect 364392 402976 364398 402988
rect 364518 402976 364524 402988
rect 364576 402976 364582 403028
rect 494054 402976 494060 403028
rect 494112 403016 494118 403028
rect 494238 403016 494244 403028
rect 494112 402988 494244 403016
rect 494112 402976 494118 402988
rect 494238 402976 494244 402988
rect 494296 402976 494302 403028
rect 299198 401548 299204 401600
rect 299256 401588 299262 401600
rect 299566 401588 299572 401600
rect 299256 401560 299572 401588
rect 299256 401548 299262 401560
rect 299566 401548 299572 401560
rect 299624 401548 299630 401600
rect 8018 398936 8024 398948
rect 7979 398908 8024 398936
rect 8018 398896 8024 398908
rect 8076 398896 8082 398948
rect 429286 398800 429292 398812
rect 429247 398772 429292 398800
rect 429286 398760 429292 398772
rect 429344 398760 429350 398812
rect 542446 398800 542452 398812
rect 542407 398772 542452 398800
rect 542446 398760 542452 398772
rect 542504 398760 542510 398812
rect 4062 394680 4068 394732
rect 4120 394720 4126 394732
rect 281626 394720 281632 394732
rect 4120 394692 281632 394720
rect 4120 394680 4126 394692
rect 281626 394680 281632 394692
rect 281684 394680 281690 394732
rect 286410 391960 286416 392012
rect 286468 392000 286474 392012
rect 580166 392000 580172 392012
rect 286468 391972 580172 392000
rect 286468 391960 286474 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 299382 391892 299388 391944
rect 299440 391932 299446 391944
rect 299569 391935 299627 391941
rect 299569 391932 299581 391935
rect 299440 391904 299581 391932
rect 299440 391892 299446 391904
rect 299569 391901 299581 391904
rect 299615 391901 299627 391935
rect 299569 391895 299627 391901
rect 8018 390572 8024 390584
rect 7979 390544 8024 390572
rect 8018 390532 8024 390544
rect 8076 390532 8082 390584
rect 429286 389172 429292 389224
rect 429344 389172 429350 389224
rect 542446 389172 542452 389224
rect 542504 389172 542510 389224
rect 429304 389088 429332 389172
rect 542464 389088 542492 389172
rect 299566 389076 299572 389088
rect 299527 389048 299572 389076
rect 299566 389036 299572 389048
rect 299624 389036 299630 389088
rect 429286 389036 429292 389088
rect 429344 389036 429350 389088
rect 542446 389036 542452 389088
rect 542504 389036 542510 389088
rect 364334 383664 364340 383716
rect 364392 383704 364398 383716
rect 364518 383704 364524 383716
rect 364392 383676 364524 383704
rect 364392 383664 364398 383676
rect 364518 383664 364524 383676
rect 364576 383664 364582 383716
rect 494054 383664 494060 383716
rect 494112 383704 494118 383716
rect 494238 383704 494244 383716
rect 494112 383676 494244 383704
rect 494112 383664 494118 383676
rect 494238 383664 494244 383676
rect 494296 383664 494302 383716
rect 7834 380876 7840 380928
rect 7892 380916 7898 380928
rect 8018 380916 8024 380928
rect 7892 380888 8024 380916
rect 7892 380876 7898 380888
rect 8018 380876 8024 380888
rect 8076 380876 8082 380928
rect 3970 379516 3976 379568
rect 4028 379556 4034 379568
rect 24118 379556 24124 379568
rect 4028 379528 24124 379556
rect 4028 379516 4034 379528
rect 24118 379516 24124 379528
rect 24176 379516 24182 379568
rect 299566 379448 299572 379500
rect 299624 379488 299630 379500
rect 299750 379488 299756 379500
rect 299624 379460 299756 379488
rect 299624 379448 299630 379460
rect 299750 379448 299756 379460
rect 299808 379448 299814 379500
rect 429286 379448 429292 379500
rect 429344 379488 429350 379500
rect 429470 379488 429476 379500
rect 429344 379460 429476 379488
rect 429344 379448 429350 379460
rect 429470 379448 429476 379460
rect 429528 379448 429534 379500
rect 542446 379448 542452 379500
rect 542504 379488 542510 379500
rect 542630 379488 542636 379500
rect 542504 379460 542636 379488
rect 542504 379448 542510 379460
rect 542630 379448 542636 379460
rect 542688 379448 542694 379500
rect 8018 369900 8024 369912
rect 7944 369872 8024 369900
rect 7944 369844 7972 369872
rect 8018 369860 8024 369872
rect 8076 369860 8082 369912
rect 7926 369792 7932 369844
rect 7984 369792 7990 369844
rect 60550 368500 60556 368552
rect 60608 368540 60614 368552
rect 580166 368540 580172 368552
rect 60608 368512 580172 368540
rect 60608 368500 60614 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 4062 365712 4068 365764
rect 4120 365752 4126 365764
rect 183554 365752 183560 365764
rect 4120 365724 183560 365752
rect 4120 365712 4126 365724
rect 183554 365712 183560 365724
rect 183612 365712 183618 365764
rect 364518 360244 364524 360256
rect 364479 360216 364524 360244
rect 364518 360204 364524 360216
rect 364576 360204 364582 360256
rect 494238 360244 494244 360256
rect 494199 360216 494244 360244
rect 494238 360204 494244 360216
rect 494296 360204 494302 360256
rect 7926 360136 7932 360188
rect 7984 360176 7990 360188
rect 8110 360176 8116 360188
rect 7984 360148 8116 360176
rect 7984 360136 7990 360148
rect 8110 360136 8116 360148
rect 8168 360136 8174 360188
rect 299842 357524 299848 357536
rect 299803 357496 299848 357524
rect 299842 357484 299848 357496
rect 299900 357484 299906 357536
rect 364518 357524 364524 357536
rect 364479 357496 364524 357524
rect 364518 357484 364524 357496
rect 364576 357484 364582 357536
rect 429562 357524 429568 357536
rect 429523 357496 429568 357524
rect 429562 357484 429568 357496
rect 429620 357484 429626 357536
rect 494238 357524 494244 357536
rect 494199 357496 494244 357524
rect 494238 357484 494244 357496
rect 494296 357484 494302 357536
rect 542722 357524 542728 357536
rect 542683 357496 542728 357524
rect 542722 357484 542728 357496
rect 542780 357484 542786 357536
rect 304350 357416 304356 357468
rect 304408 357456 304414 357468
rect 580166 357456 580172 357468
rect 304408 357428 580172 357456
rect 304408 357416 304414 357428
rect 580166 357416 580172 357428
rect 580224 357416 580230 357468
rect 8021 357391 8079 357397
rect 8021 357357 8033 357391
rect 8067 357388 8079 357391
rect 8110 357388 8116 357400
rect 8067 357360 8116 357388
rect 8067 357357 8079 357360
rect 8021 357351 8079 357357
rect 8110 357348 8116 357360
rect 8168 357348 8174 357400
rect 299750 356124 299756 356176
rect 299808 356164 299814 356176
rect 299845 356167 299903 356173
rect 299845 356164 299857 356167
rect 299808 356136 299857 356164
rect 299808 356124 299814 356136
rect 299845 356133 299857 356136
rect 299891 356133 299903 356167
rect 299845 356127 299903 356133
rect 299842 354668 299848 354680
rect 299803 354640 299848 354668
rect 299842 354628 299848 354640
rect 299900 354628 299906 354680
rect 429562 353376 429568 353388
rect 429523 353348 429568 353376
rect 429562 353336 429568 353348
rect 429620 353336 429626 353388
rect 542722 353376 542728 353388
rect 542683 353348 542728 353376
rect 542722 353336 542728 353348
rect 542780 353336 542786 353388
rect 429654 353240 429660 353252
rect 429615 353212 429660 353240
rect 429654 353200 429660 353212
rect 429712 353200 429718 353252
rect 542814 353240 542820 353252
rect 542775 353212 542820 353240
rect 542814 353200 542820 353212
rect 542872 353200 542878 353252
rect 8018 347800 8024 347812
rect 7979 347772 8024 347800
rect 8018 347760 8024 347772
rect 8076 347760 8082 347812
rect 364334 347732 364340 347744
rect 364295 347704 364340 347732
rect 364334 347692 364340 347704
rect 364392 347692 364398 347744
rect 494054 347732 494060 347744
rect 494015 347704 494060 347732
rect 494054 347692 494060 347704
rect 494112 347692 494118 347744
rect 285122 345040 285128 345092
rect 285180 345080 285186 345092
rect 580166 345080 580172 345092
rect 285180 345052 580172 345080
rect 285180 345040 285186 345052
rect 580166 345040 580172 345052
rect 580224 345040 580230 345092
rect 8018 341000 8024 341012
rect 7979 340972 8024 341000
rect 8018 340960 8024 340972
rect 8076 340960 8082 341012
rect 429654 340796 429660 340808
rect 429615 340768 429660 340796
rect 429654 340756 429660 340768
rect 429712 340756 429718 340808
rect 542814 340796 542820 340808
rect 542775 340768 542820 340796
rect 542814 340756 542820 340768
rect 542872 340756 542878 340808
rect 364337 338147 364395 338153
rect 364337 338113 364349 338147
rect 364383 338144 364395 338147
rect 364426 338144 364432 338156
rect 364383 338116 364432 338144
rect 364383 338113 364395 338116
rect 364337 338107 364395 338113
rect 364426 338104 364432 338116
rect 364484 338104 364490 338156
rect 494057 338147 494115 338153
rect 494057 338113 494069 338147
rect 494103 338144 494115 338147
rect 494146 338144 494152 338156
rect 494103 338116 494152 338144
rect 494103 338113 494115 338116
rect 494057 338107 494115 338113
rect 494146 338104 494152 338116
rect 494204 338104 494210 338156
rect 8018 336852 8024 336864
rect 7979 336824 8024 336852
rect 8018 336812 8024 336824
rect 8076 336812 8082 336864
rect 4062 336744 4068 336796
rect 4120 336784 4126 336796
rect 281902 336784 281908 336796
rect 4120 336756 281908 336784
rect 4120 336744 4126 336756
rect 281902 336744 281908 336756
rect 281960 336744 281966 336796
rect 299845 336787 299903 336793
rect 299845 336753 299857 336787
rect 299891 336784 299903 336787
rect 299934 336784 299940 336796
rect 299891 336756 299940 336784
rect 299891 336753 299903 336756
rect 299845 336747 299903 336753
rect 299934 336744 299940 336756
rect 299992 336744 299998 336796
rect 7929 336651 7987 336657
rect 7929 336617 7941 336651
rect 7975 336648 7987 336651
rect 8018 336648 8024 336660
rect 7975 336620 8024 336648
rect 7975 336617 7987 336620
rect 7929 336611 7987 336617
rect 8018 336608 8024 336620
rect 8076 336608 8082 336660
rect 7926 327128 7932 327140
rect 7887 327100 7932 327128
rect 7926 327088 7932 327100
rect 7984 327088 7990 327140
rect 299750 327088 299756 327140
rect 299808 327128 299814 327140
rect 299842 327128 299848 327140
rect 299808 327100 299848 327128
rect 299808 327088 299814 327100
rect 299842 327088 299848 327100
rect 299900 327088 299906 327140
rect 364334 325660 364340 325712
rect 364392 325700 364398 325712
rect 364518 325700 364524 325712
rect 364392 325672 364524 325700
rect 364392 325660 364398 325672
rect 364518 325660 364524 325672
rect 364576 325660 364582 325712
rect 429470 325660 429476 325712
rect 429528 325700 429534 325712
rect 429562 325700 429568 325712
rect 429528 325672 429568 325700
rect 429528 325660 429534 325672
rect 429562 325660 429568 325672
rect 429620 325660 429626 325712
rect 494054 325660 494060 325712
rect 494112 325700 494118 325712
rect 494238 325700 494244 325712
rect 494112 325672 494244 325700
rect 494112 325660 494118 325672
rect 494238 325660 494244 325672
rect 494296 325660 494302 325712
rect 542630 325660 542636 325712
rect 542688 325700 542694 325712
rect 542722 325700 542728 325712
rect 542688 325672 542728 325700
rect 542688 325660 542694 325672
rect 542722 325660 542728 325672
rect 542780 325660 542786 325712
rect 291930 321580 291936 321632
rect 291988 321620 291994 321632
rect 580166 321620 580172 321632
rect 291988 321592 580172 321620
rect 291988 321580 291994 321592
rect 580166 321580 580172 321592
rect 580224 321580 580230 321632
rect 7926 321444 7932 321496
rect 7984 321484 7990 321496
rect 8202 321484 8208 321496
rect 7984 321456 8208 321484
rect 7984 321444 7990 321456
rect 8202 321444 8208 321456
rect 8260 321444 8266 321496
rect 299658 318792 299664 318844
rect 299716 318832 299722 318844
rect 299750 318832 299756 318844
rect 299716 318804 299756 318832
rect 299716 318792 299722 318804
rect 299750 318792 299756 318804
rect 299808 318792 299814 318844
rect 429378 318792 429384 318844
rect 429436 318832 429442 318844
rect 429470 318832 429476 318844
rect 429436 318804 429476 318832
rect 429436 318792 429442 318804
rect 429470 318792 429476 318804
rect 429528 318792 429534 318844
rect 542538 318792 542544 318844
rect 542596 318832 542602 318844
rect 542630 318832 542636 318844
rect 542596 318804 542636 318832
rect 542596 318792 542602 318804
rect 542630 318792 542636 318804
rect 542688 318792 542694 318844
rect 299658 311924 299664 311976
rect 299716 311964 299722 311976
rect 299750 311964 299756 311976
rect 299716 311936 299756 311964
rect 299716 311924 299722 311936
rect 299750 311924 299756 311936
rect 299808 311924 299814 311976
rect 429378 311924 429384 311976
rect 429436 311964 429442 311976
rect 429470 311964 429476 311976
rect 429436 311936 429476 311964
rect 429436 311924 429442 311936
rect 429470 311924 429476 311936
rect 429528 311924 429534 311976
rect 542538 311924 542544 311976
rect 542596 311964 542602 311976
rect 542630 311964 542636 311976
rect 542596 311936 542636 311964
rect 542596 311924 542602 311936
rect 542630 311924 542636 311936
rect 542688 311924 542694 311976
rect 61194 310496 61200 310548
rect 61252 310536 61258 310548
rect 579798 310536 579804 310548
rect 61252 310508 579804 310536
rect 61252 310496 61258 310508
rect 579798 310496 579804 310508
rect 579856 310496 579862 310548
rect 7926 309204 7932 309256
rect 7984 309244 7990 309256
rect 8202 309244 8208 309256
rect 7984 309216 8208 309244
rect 7984 309204 7990 309216
rect 8202 309204 8208 309216
rect 8260 309204 8266 309256
rect 4062 307776 4068 307828
rect 4120 307816 4126 307828
rect 22738 307816 22744 307828
rect 4120 307788 22744 307816
rect 4120 307776 4126 307788
rect 22738 307776 22744 307788
rect 22796 307776 22802 307828
rect 364334 306348 364340 306400
rect 364392 306388 364398 306400
rect 364518 306388 364524 306400
rect 364392 306360 364524 306388
rect 364392 306348 364398 306360
rect 364518 306348 364524 306360
rect 364576 306348 364582 306400
rect 494054 306348 494060 306400
rect 494112 306388 494118 306400
rect 494238 306388 494244 306400
rect 494112 306360 494244 306388
rect 494112 306348 494118 306360
rect 494238 306348 494244 306360
rect 494296 306348 494302 306400
rect 8018 302268 8024 302320
rect 8076 302268 8082 302320
rect 8036 302104 8064 302268
rect 299566 302200 299572 302252
rect 299624 302240 299630 302252
rect 299750 302240 299756 302252
rect 299624 302212 299756 302240
rect 299624 302200 299630 302212
rect 299750 302200 299756 302212
rect 299808 302200 299814 302252
rect 429286 302200 429292 302252
rect 429344 302240 429350 302252
rect 429470 302240 429476 302252
rect 429344 302212 429476 302240
rect 429344 302200 429350 302212
rect 429470 302200 429476 302212
rect 429528 302200 429534 302252
rect 542446 302200 542452 302252
rect 542504 302240 542510 302252
rect 542630 302240 542636 302252
rect 542504 302212 542636 302240
rect 542504 302200 542510 302212
rect 542630 302200 542636 302212
rect 542688 302200 542694 302252
rect 8110 302104 8116 302116
rect 8036 302076 8116 302104
rect 8110 302064 8116 302076
rect 8168 302064 8174 302116
rect 299658 299452 299664 299464
rect 299619 299424 299664 299452
rect 299658 299412 299664 299424
rect 299716 299412 299722 299464
rect 216582 298120 216588 298172
rect 216640 298160 216646 298172
rect 580166 298160 580172 298172
rect 216640 298132 580172 298160
rect 216640 298120 216646 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3142 293972 3148 294024
rect 3200 294012 3206 294024
rect 7558 294012 7564 294024
rect 3200 293984 7564 294012
rect 3200 293972 3206 293984
rect 7558 293972 7564 293984
rect 7616 293972 7622 294024
rect 299661 289867 299719 289873
rect 299661 289833 299673 289867
rect 299707 289864 299719 289867
rect 299750 289864 299756 289876
rect 299707 289836 299756 289864
rect 299707 289833 299719 289836
rect 299661 289827 299719 289833
rect 299750 289824 299756 289836
rect 299808 289824 299814 289876
rect 8113 289799 8171 289805
rect 8113 289765 8125 289799
rect 8159 289796 8171 289799
rect 8202 289796 8208 289808
rect 8159 289768 8208 289796
rect 8159 289765 8171 289768
rect 8113 289759 8171 289765
rect 8202 289756 8208 289768
rect 8260 289756 8266 289808
rect 429470 289796 429476 289808
rect 429431 289768 429476 289796
rect 429470 289756 429476 289768
rect 429528 289756 429534 289808
rect 542449 289799 542507 289805
rect 542449 289765 542461 289799
rect 542495 289796 542507 289799
rect 542630 289796 542636 289808
rect 542495 289768 542636 289796
rect 542495 289765 542507 289768
rect 542449 289759 542507 289765
rect 542630 289756 542636 289768
rect 542688 289756 542694 289808
rect 364334 287036 364340 287088
rect 364392 287076 364398 287088
rect 364518 287076 364524 287088
rect 364392 287048 364524 287076
rect 364392 287036 364398 287048
rect 364518 287036 364524 287048
rect 364576 287036 364582 287088
rect 494054 287036 494060 287088
rect 494112 287076 494118 287088
rect 494238 287076 494244 287088
rect 494112 287048 494244 287076
rect 494112 287036 494118 287048
rect 494238 287036 494244 287048
rect 494296 287036 494302 287088
rect 286502 282140 286508 282192
rect 286560 282180 286566 282192
rect 494054 282180 494060 282192
rect 286560 282152 494060 282180
rect 286560 282140 286566 282152
rect 494054 282140 494060 282152
rect 494112 282140 494118 282192
rect 8110 280208 8116 280220
rect 8071 280180 8116 280208
rect 8110 280168 8116 280180
rect 8168 280168 8174 280220
rect 429473 280211 429531 280217
rect 429473 280177 429485 280211
rect 429519 280208 429531 280211
rect 429562 280208 429568 280220
rect 429519 280180 429568 280208
rect 429519 280177 429531 280180
rect 429473 280171 429531 280177
rect 429562 280168 429568 280180
rect 429620 280168 429626 280220
rect 542446 280208 542452 280220
rect 542407 280180 542452 280208
rect 542446 280168 542452 280180
rect 542504 280168 542510 280220
rect 89622 277992 89628 278044
rect 89680 278032 89686 278044
rect 283374 278032 283380 278044
rect 89680 278004 283380 278032
rect 89680 277992 89686 278004
rect 283374 277992 283380 278004
rect 283432 277992 283438 278044
rect 429378 274864 429384 274916
rect 429436 274904 429442 274916
rect 429562 274904 429568 274916
rect 429436 274876 429568 274904
rect 429436 274864 429442 274876
rect 429562 274864 429568 274876
rect 429620 274864 429626 274916
rect 290550 274660 290556 274712
rect 290608 274700 290614 274712
rect 580166 274700 580172 274712
rect 290608 274672 580172 274700
rect 290608 274660 290614 274672
rect 580166 274660 580172 274672
rect 580224 274660 580230 274712
rect 202782 273912 202788 273964
rect 202840 273952 202846 273964
rect 283466 273952 283472 273964
rect 202840 273924 283472 273952
rect 202840 273912 202846 273924
rect 283466 273912 283472 273924
rect 283524 273912 283530 273964
rect 8110 273300 8116 273352
rect 8168 273300 8174 273352
rect 8128 273148 8156 273300
rect 8110 273096 8116 273148
rect 8168 273096 8174 273148
rect 60458 272484 60464 272536
rect 60516 272524 60522 272536
rect 462314 272524 462320 272536
rect 60516 272496 462320 272524
rect 60516 272484 60522 272496
rect 462314 272484 462320 272496
rect 462372 272484 462378 272536
rect 60918 271124 60924 271176
rect 60976 271164 60982 271176
rect 527174 271164 527180 271176
rect 60976 271136 527180 271164
rect 60976 271124 60982 271136
rect 527174 271124 527180 271136
rect 527232 271124 527238 271176
rect 98638 270648 98644 270700
rect 98696 270688 98702 270700
rect 442994 270688 443000 270700
rect 98696 270660 443000 270688
rect 98696 270648 98702 270660
rect 442994 270648 443000 270660
rect 443052 270648 443058 270700
rect 64046 270580 64052 270632
rect 64104 270620 64110 270632
rect 458174 270620 458180 270632
rect 64104 270592 458180 270620
rect 64104 270580 64110 270592
rect 458174 270580 458180 270592
rect 458232 270580 458238 270632
rect 73798 270512 73804 270564
rect 73856 270552 73862 270564
rect 476114 270552 476120 270564
rect 73856 270524 476120 270552
rect 73856 270512 73862 270524
rect 476114 270512 476120 270524
rect 476172 270512 476178 270564
rect 429378 270484 429384 270496
rect 429339 270456 429384 270484
rect 429378 270444 429384 270456
rect 429436 270444 429442 270496
rect 97534 269968 97540 270020
rect 97592 270008 97598 270020
rect 460934 270008 460940 270020
rect 97592 269980 460940 270008
rect 97592 269968 97598 269980
rect 460934 269968 460940 269980
rect 460992 269968 460998 270020
rect 120350 269900 120356 269952
rect 120408 269940 120414 269952
rect 520274 269940 520280 269952
rect 120408 269912 520280 269940
rect 120408 269900 120414 269912
rect 520274 269900 520280 269912
rect 520332 269900 520338 269952
rect 189534 269832 189540 269884
rect 189592 269872 189598 269884
rect 285950 269872 285956 269884
rect 189592 269844 285956 269872
rect 189592 269832 189598 269844
rect 285950 269832 285956 269844
rect 286008 269832 286014 269884
rect 22738 269764 22744 269816
rect 22796 269804 22802 269816
rect 76742 269804 76748 269816
rect 22796 269776 76748 269804
rect 22796 269764 22802 269776
rect 76742 269764 76748 269776
rect 76800 269764 76806 269816
rect 187694 269764 187700 269816
rect 187752 269804 187758 269816
rect 289814 269804 289820 269816
rect 187752 269776 289820 269804
rect 187752 269764 187758 269776
rect 289814 269764 289820 269776
rect 289872 269764 289878 269816
rect 164878 269696 164884 269748
rect 164936 269736 164942 269748
rect 288526 269736 288532 269748
rect 164936 269708 288532 269736
rect 164936 269696 164942 269708
rect 288526 269696 288532 269708
rect 288584 269696 288590 269748
rect 156966 269628 156972 269680
rect 157024 269668 157030 269680
rect 287146 269668 287152 269680
rect 157024 269640 287152 269668
rect 157024 269628 157030 269640
rect 287146 269628 287152 269640
rect 287204 269628 287210 269680
rect 152918 269560 152924 269612
rect 152976 269600 152982 269612
rect 285674 269600 285680 269612
rect 152976 269572 285680 269600
rect 152976 269560 152982 269572
rect 285674 269560 285680 269572
rect 285732 269560 285738 269612
rect 181622 269492 181628 269544
rect 181680 269532 181686 269544
rect 412634 269532 412640 269544
rect 181680 269504 412640 269532
rect 181680 269492 181686 269504
rect 412634 269492 412640 269504
rect 412692 269492 412698 269544
rect 174814 269424 174820 269476
rect 174872 269464 174878 269476
rect 418154 269464 418160 269476
rect 174872 269436 418160 269464
rect 174872 269424 174878 269436
rect 418154 269424 418160 269436
rect 418212 269424 418218 269476
rect 139118 269356 139124 269408
rect 139176 269396 139182 269408
rect 416866 269396 416872 269408
rect 139176 269368 416872 269396
rect 139176 269356 139182 269368
rect 416866 269356 416872 269368
rect 416924 269356 416930 269408
rect 163958 269288 163964 269340
rect 164016 269328 164022 269340
rect 465074 269328 465080 269340
rect 164016 269300 465080 269328
rect 164016 269288 164022 269300
rect 465074 269288 465080 269300
rect 465132 269288 465138 269340
rect 112438 269220 112444 269272
rect 112496 269260 112502 269272
rect 419534 269260 419540 269272
rect 112496 269232 419540 269260
rect 112496 269220 112502 269232
rect 419534 269220 419540 269232
rect 419592 269220 419598 269272
rect 262766 269152 262772 269204
rect 262824 269192 262830 269204
rect 287238 269192 287244 269204
rect 262824 269164 287244 269192
rect 262824 269152 262830 269164
rect 287238 269152 287244 269164
rect 287296 269152 287302 269204
rect 260742 269084 260748 269136
rect 260800 269124 260806 269136
rect 286042 269124 286048 269136
rect 260800 269096 286048 269124
rect 260800 269084 260806 269096
rect 286042 269084 286048 269096
rect 286100 269084 286106 269136
rect 163038 268608 163044 268660
rect 163096 268648 163102 268660
rect 542446 268648 542452 268660
rect 163096 268620 542452 268648
rect 163096 268608 163102 268620
rect 542446 268608 542452 268620
rect 542504 268608 542510 268660
rect 220262 268540 220268 268592
rect 220320 268580 220326 268592
rect 294690 268580 294696 268592
rect 220320 268552 294696 268580
rect 220320 268540 220326 268552
rect 294690 268540 294696 268552
rect 294748 268540 294754 268592
rect 211430 268472 211436 268524
rect 211488 268512 211494 268524
rect 293310 268512 293316 268524
rect 211488 268484 293316 268512
rect 211488 268472 211494 268484
rect 293310 268472 293316 268484
rect 293368 268472 293374 268524
rect 172790 268404 172796 268456
rect 172848 268444 172854 268456
rect 281810 268444 281816 268456
rect 172848 268416 281816 268444
rect 172848 268404 172854 268416
rect 281810 268404 281816 268416
rect 281868 268404 281874 268456
rect 178678 268336 178684 268388
rect 178736 268376 178742 268388
rect 288618 268376 288624 268388
rect 178736 268348 288624 268376
rect 178736 268336 178742 268348
rect 288618 268336 288624 268348
rect 288676 268336 288682 268388
rect 213270 268268 213276 268320
rect 213328 268308 213334 268320
rect 408494 268308 408500 268320
rect 213328 268280 408500 268308
rect 213328 268268 213334 268280
rect 408494 268268 408500 268280
rect 408552 268268 408558 268320
rect 55858 268200 55864 268252
rect 55916 268240 55922 268252
rect 214374 268240 214380 268252
rect 55916 268212 214380 268240
rect 55916 268200 55922 268212
rect 214374 268200 214380 268212
rect 214432 268200 214438 268252
rect 236086 268200 236092 268252
rect 236144 268240 236150 268252
rect 436094 268240 436100 268252
rect 236144 268212 436100 268240
rect 236144 268200 236150 268212
rect 436094 268200 436100 268212
rect 436152 268200 436158 268252
rect 69014 268132 69020 268184
rect 69072 268172 69078 268184
rect 283282 268172 283288 268184
rect 69072 268144 283288 268172
rect 69072 268132 69078 268144
rect 283282 268132 283288 268144
rect 283340 268132 283346 268184
rect 6270 268064 6276 268116
rect 6328 268104 6334 268116
rect 273622 268104 273628 268116
rect 6328 268076 273628 268104
rect 6328 268064 6334 268076
rect 273622 268064 273628 268076
rect 273680 268064 273686 268116
rect 168742 267996 168748 268048
rect 168800 268036 168806 268048
rect 518894 268036 518900 268048
rect 168800 268008 518900 268036
rect 168800 267996 168806 268008
rect 518894 267996 518900 268008
rect 518952 267996 518958 268048
rect 19978 267928 19984 267980
rect 20036 267968 20042 267980
rect 229094 267968 229100 267980
rect 20036 267940 229100 267968
rect 20036 267928 20042 267940
rect 229094 267928 229100 267940
rect 229152 267928 229158 267980
rect 230198 267928 230204 267980
rect 230256 267968 230262 267980
rect 579798 267968 579804 267980
rect 230256 267940 579804 267968
rect 230256 267928 230262 267940
rect 579798 267928 579804 267940
rect 579856 267928 579862 267980
rect 188614 267860 188620 267912
rect 188672 267900 188678 267912
rect 539594 267900 539600 267912
rect 188672 267872 539600 267900
rect 188672 267860 188678 267872
rect 539594 267860 539600 267872
rect 539652 267860 539658 267912
rect 145006 267792 145012 267844
rect 145064 267832 145070 267844
rect 521654 267832 521660 267844
rect 145064 267804 521660 267832
rect 145064 267792 145070 267804
rect 521654 267792 521660 267804
rect 521712 267792 521718 267844
rect 252830 267724 252836 267776
rect 252888 267764 252894 267776
rect 284386 267764 284392 267776
rect 252888 267736 284392 267764
rect 252888 267724 252894 267736
rect 284386 267724 284392 267736
rect 284444 267724 284450 267776
rect 542354 267724 542360 267776
rect 542412 267764 542418 267776
rect 542630 267764 542636 267776
rect 542412 267736 542636 267764
rect 542412 267724 542418 267736
rect 542630 267724 542636 267736
rect 542688 267724 542694 267776
rect 99558 267656 99564 267708
rect 99616 267696 99622 267708
rect 100662 267696 100668 267708
rect 99616 267668 100668 267696
rect 99616 267656 99622 267668
rect 100662 267656 100668 267668
rect 100720 267656 100726 267708
rect 110414 267656 110420 267708
rect 110472 267696 110478 267708
rect 111702 267696 111708 267708
rect 110472 267668 111708 267696
rect 110472 267656 110478 267668
rect 111702 267656 111708 267668
rect 111760 267656 111766 267708
rect 248966 267656 248972 267708
rect 249024 267696 249030 267708
rect 249702 267696 249708 267708
rect 249024 267668 249708 267696
rect 249024 267656 249030 267668
rect 249702 267656 249708 267668
rect 249760 267656 249766 267708
rect 280614 267656 280620 267708
rect 280672 267696 280678 267708
rect 281442 267696 281448 267708
rect 280672 267668 281448 267696
rect 280672 267656 280678 267668
rect 281442 267656 281448 267668
rect 281500 267656 281506 267708
rect 89622 267316 89628 267368
rect 89680 267356 89686 267368
rect 270494 267356 270500 267368
rect 89680 267328 270500 267356
rect 89680 267316 89686 267328
rect 270494 267316 270500 267328
rect 270552 267316 270558 267368
rect 259822 267248 259828 267300
rect 259880 267288 259886 267300
rect 281350 267288 281356 267300
rect 259880 267260 281356 267288
rect 259880 267248 259886 267260
rect 281350 267248 281356 267260
rect 281408 267248 281414 267300
rect 115382 267180 115388 267232
rect 115440 267220 115446 267232
rect 257982 267220 257988 267232
rect 115440 267192 257988 267220
rect 115440 267180 115446 267192
rect 257982 267180 257988 267192
rect 258040 267180 258046 267232
rect 263686 267180 263692 267232
rect 263744 267220 263750 267232
rect 287882 267220 287888 267232
rect 263744 267192 287888 267220
rect 263744 267180 263750 267192
rect 287882 267180 287888 267192
rect 287940 267180 287946 267232
rect 249886 267112 249892 267164
rect 249944 267152 249950 267164
rect 282270 267152 282276 267164
rect 249944 267124 282276 267152
rect 249944 267112 249950 267124
rect 282270 267112 282276 267124
rect 282328 267112 282334 267164
rect 84654 267044 84660 267096
rect 84712 267084 84718 267096
rect 304994 267084 305000 267096
rect 84712 267056 305000 267084
rect 84712 267044 84718 267056
rect 304994 267044 305000 267056
rect 305052 267044 305058 267096
rect 57698 266976 57704 267028
rect 57756 267016 57762 267028
rect 116302 267016 116308 267028
rect 57756 266988 116308 267016
rect 57756 266976 57762 266988
rect 116302 266976 116308 266988
rect 116360 266976 116366 267028
rect 265710 266976 265716 267028
rect 265768 267016 265774 267028
rect 281166 267016 281172 267028
rect 265768 266988 281172 267016
rect 265768 266976 265774 266988
rect 281166 266976 281172 266988
rect 281224 266976 281230 267028
rect 57790 266908 57796 266960
rect 57848 266948 57854 266960
rect 128262 266948 128268 266960
rect 57848 266920 128268 266948
rect 57848 266908 57854 266920
rect 128262 266908 128268 266920
rect 128320 266908 128326 266960
rect 132862 266908 132868 266960
rect 132920 266948 132926 266960
rect 180702 266948 180708 266960
rect 132920 266920 180708 266948
rect 132920 266908 132926 266920
rect 180702 266908 180708 266920
rect 180760 266908 180766 266960
rect 237006 266908 237012 266960
rect 237064 266948 237070 266960
rect 281718 266948 281724 266960
rect 237064 266920 281724 266948
rect 237064 266908 237070 266920
rect 281718 266908 281724 266920
rect 281776 266908 281782 266960
rect 57882 266840 57888 266892
rect 57940 266880 57946 266892
rect 137094 266880 137100 266892
rect 57940 266852 137100 266880
rect 57940 266840 57946 266852
rect 137094 266840 137100 266852
rect 137152 266840 137158 266892
rect 226150 266840 226156 266892
rect 226208 266880 226214 266892
rect 287790 266880 287796 266892
rect 226208 266852 287796 266880
rect 226208 266840 226214 266852
rect 287790 266840 287796 266852
rect 287848 266840 287854 266892
rect 56318 266772 56324 266824
rect 56376 266812 56382 266824
rect 154942 266812 154948 266824
rect 56376 266784 154948 266812
rect 56376 266772 56382 266784
rect 154942 266772 154948 266784
rect 155000 266772 155006 266824
rect 164142 266772 164148 266824
rect 164200 266812 164206 266824
rect 197446 266812 197452 266824
rect 164200 266784 197452 266812
rect 164200 266772 164206 266784
rect 197446 266772 197452 266784
rect 197504 266772 197510 266824
rect 198550 266772 198556 266824
rect 198608 266812 198614 266824
rect 281994 266812 282000 266824
rect 198608 266784 282000 266812
rect 198608 266772 198614 266784
rect 281994 266772 282000 266784
rect 282052 266772 282058 266824
rect 56226 266704 56232 266756
rect 56284 266744 56290 266756
rect 179782 266744 179788 266756
rect 56284 266716 179788 266744
rect 56284 266704 56290 266716
rect 179782 266704 179788 266716
rect 179840 266704 179846 266756
rect 194502 266704 194508 266756
rect 194560 266744 194566 266756
rect 282454 266744 282460 266756
rect 194560 266716 282460 266744
rect 194560 266704 194566 266716
rect 282454 266704 282460 266716
rect 282512 266704 282518 266756
rect 67910 266636 67916 266688
rect 67968 266676 67974 266688
rect 126974 266676 126980 266688
rect 67968 266648 126980 266676
rect 67968 266636 67974 266648
rect 126974 266636 126980 266648
rect 127032 266636 127038 266688
rect 256878 266636 256884 266688
rect 256936 266676 256942 266688
rect 283098 266676 283104 266688
rect 256936 266648 283104 266676
rect 256936 266636 256942 266648
rect 283098 266636 283104 266648
rect 283156 266636 283162 266688
rect 17218 266568 17224 266620
rect 17276 266608 17282 266620
rect 117406 266608 117412 266620
rect 17276 266580 117412 266608
rect 17276 266568 17282 266580
rect 117406 266568 117412 266580
rect 117464 266568 117470 266620
rect 124214 266568 124220 266620
rect 124272 266608 124278 266620
rect 282362 266608 282368 266620
rect 124272 266580 282368 266608
rect 124272 266568 124278 266580
rect 282362 266568 282368 266580
rect 282420 266568 282426 266620
rect 157886 266500 157892 266552
rect 157944 266540 157950 266552
rect 160097 266543 160155 266549
rect 160097 266540 160109 266543
rect 157944 266512 160109 266540
rect 157944 266500 157950 266512
rect 160097 266509 160109 266512
rect 160143 266509 160155 266543
rect 160097 266503 160155 266509
rect 270678 266500 270684 266552
rect 270736 266540 270742 266552
rect 283558 266540 283564 266552
rect 270736 266512 283564 266540
rect 270736 266500 270742 266512
rect 283558 266500 283564 266512
rect 283616 266500 283622 266552
rect 55122 266432 55128 266484
rect 55180 266472 55186 266484
rect 66990 266472 66996 266484
rect 55180 266444 66996 266472
rect 55180 266432 55186 266444
rect 66990 266432 66996 266444
rect 67048 266432 67054 266484
rect 71958 266432 71964 266484
rect 72016 266472 72022 266484
rect 259454 266472 259460 266484
rect 72016 266444 259460 266472
rect 72016 266432 72022 266444
rect 259454 266432 259460 266444
rect 259512 266432 259518 266484
rect 267734 266432 267740 266484
rect 267792 266472 267798 266484
rect 288710 266472 288716 266484
rect 267792 266444 288716 266472
rect 267792 266432 267798 266444
rect 288710 266432 288716 266444
rect 288768 266432 288774 266484
rect 53742 266364 53748 266416
rect 53800 266404 53806 266416
rect 65886 266404 65892 266416
rect 53800 266376 65892 266404
rect 53800 266364 53806 266376
rect 65886 266364 65892 266376
rect 65944 266364 65950 266416
rect 122374 266364 122380 266416
rect 122432 266404 122438 266416
rect 128354 266404 128360 266416
rect 122432 266376 128360 266404
rect 122432 266364 122438 266376
rect 128354 266364 128360 266376
rect 128412 266364 128418 266416
rect 158990 266364 158996 266416
rect 159048 266404 159054 266416
rect 160002 266404 160008 266416
rect 159048 266376 160008 266404
rect 159048 266364 159054 266376
rect 160002 266364 160008 266376
rect 160060 266364 160066 266416
rect 160097 266407 160155 266413
rect 160097 266373 160109 266407
rect 160143 266404 160155 266407
rect 163406 266404 163412 266416
rect 160143 266376 163412 266404
rect 160143 266373 160155 266376
rect 160097 266367 160155 266373
rect 163406 266364 163412 266376
rect 163464 266364 163470 266416
rect 210326 266364 210332 266416
rect 210384 266404 210390 266416
rect 226242 266404 226248 266416
rect 210384 266376 226248 266404
rect 210384 266364 210390 266376
rect 226242 266364 226248 266376
rect 226300 266364 226306 266416
rect 277670 266364 277676 266416
rect 277728 266404 277734 266416
rect 280890 266404 280896 266416
rect 277728 266376 280896 266404
rect 277728 266364 277734 266376
rect 280890 266364 280896 266376
rect 280948 266364 280954 266416
rect 3878 266296 3884 266348
rect 3936 266336 3942 266348
rect 69014 266336 69020 266348
rect 3936 266308 69020 266336
rect 3936 266296 3942 266308
rect 69014 266296 69020 266308
rect 69072 266296 69078 266348
rect 263594 266296 263600 266348
rect 263652 266336 263658 266348
rect 263652 266308 263697 266336
rect 263652 266296 263658 266308
rect 271782 266268 271788 266280
rect 271743 266240 271788 266268
rect 271782 266228 271788 266240
rect 271840 266228 271846 266280
rect 155862 265820 155868 265872
rect 155920 265860 155926 265872
rect 482278 265860 482284 265872
rect 155920 265832 482284 265860
rect 155920 265820 155926 265832
rect 482278 265820 482284 265832
rect 482336 265820 482342 265872
rect 231118 265752 231124 265804
rect 231176 265792 231182 265804
rect 284294 265792 284300 265804
rect 231176 265764 284300 265792
rect 231176 265752 231182 265764
rect 284294 265752 284300 265764
rect 284352 265752 284358 265804
rect 3510 265684 3516 265736
rect 3568 265724 3574 265736
rect 164142 265724 164148 265736
rect 3568 265696 164148 265724
rect 3568 265684 3574 265696
rect 164142 265684 164148 265696
rect 164200 265684 164206 265736
rect 257982 265684 257988 265736
rect 258040 265724 258046 265736
rect 373994 265724 374000 265736
rect 258040 265696 374000 265724
rect 258040 265684 258046 265696
rect 373994 265684 374000 265696
rect 374052 265684 374058 265736
rect 128354 265616 128360 265668
rect 128412 265656 128418 265668
rect 351914 265656 351920 265668
rect 128412 265628 351920 265656
rect 128412 265616 128418 265628
rect 351914 265616 351920 265628
rect 351972 265616 351978 265668
rect 275646 265548 275652 265600
rect 275704 265588 275710 265600
rect 345014 265588 345020 265600
rect 275704 265560 345020 265588
rect 275704 265548 275710 265560
rect 345014 265548 345020 265560
rect 345072 265548 345078 265600
rect 215294 265480 215300 265532
rect 215352 265520 215358 265532
rect 286134 265520 286140 265532
rect 215352 265492 286140 265520
rect 215352 265480 215358 265492
rect 286134 265480 286140 265492
rect 286192 265480 286198 265532
rect 221182 265412 221188 265464
rect 221240 265452 221246 265464
rect 298094 265452 298100 265464
rect 221240 265424 298100 265452
rect 221240 265412 221246 265424
rect 298094 265412 298100 265424
rect 298152 265412 298158 265464
rect 149974 265344 149980 265396
rect 150032 265384 150038 265396
rect 284570 265384 284576 265396
rect 150032 265356 284576 265384
rect 150032 265344 150038 265356
rect 284570 265344 284576 265356
rect 284628 265344 284634 265396
rect 96614 265276 96620 265328
rect 96672 265316 96678 265328
rect 327074 265316 327080 265328
rect 96672 265288 327080 265316
rect 96672 265276 96678 265288
rect 327074 265276 327080 265288
rect 327132 265276 327138 265328
rect 171870 265208 171876 265260
rect 171928 265248 171934 265260
rect 437474 265248 437480 265260
rect 171928 265220 437480 265248
rect 171928 265208 171934 265220
rect 437474 265208 437480 265220
rect 437532 265208 437538 265260
rect 161934 265140 161940 265192
rect 161992 265180 161998 265192
rect 435358 265180 435364 265192
rect 161992 265152 435364 265180
rect 161992 265140 161998 265152
rect 435358 265140 435364 265152
rect 435416 265140 435422 265192
rect 68830 265072 68836 265124
rect 68888 265112 68894 265124
rect 347774 265112 347780 265124
rect 68888 265084 347780 265112
rect 68888 265072 68894 265084
rect 347774 265072 347780 265084
rect 347832 265072 347838 265124
rect 233050 265004 233056 265056
rect 233108 265044 233114 265056
rect 547874 265044 547880 265056
rect 233108 265016 547880 265044
rect 233108 265004 233114 265016
rect 547874 265004 547880 265016
rect 547932 265004 547938 265056
rect 268930 264936 268936 264988
rect 268988 264976 268994 264988
rect 287054 264976 287060 264988
rect 268988 264948 287060 264976
rect 268988 264936 268994 264948
rect 287054 264936 287060 264948
rect 287112 264936 287118 264988
rect 277949 264639 278007 264645
rect 277949 264605 277961 264639
rect 277995 264636 278007 264639
rect 285766 264636 285772 264648
rect 277995 264608 285772 264636
rect 277995 264605 278007 264608
rect 277949 264599 278007 264605
rect 285766 264596 285772 264608
rect 285824 264596 285830 264648
rect 9677 264571 9735 264577
rect 9677 264537 9689 264571
rect 9723 264568 9735 264571
rect 19245 264571 19303 264577
rect 19245 264568 19257 264571
rect 9723 264540 19257 264568
rect 9723 264537 9735 264540
rect 9677 264531 9735 264537
rect 19245 264537 19257 264540
rect 19291 264537 19303 264571
rect 19245 264531 19303 264537
rect 28997 264571 29055 264577
rect 28997 264537 29009 264571
rect 29043 264568 29055 264571
rect 38565 264571 38623 264577
rect 38565 264568 38577 264571
rect 29043 264540 38577 264568
rect 29043 264537 29055 264540
rect 28997 264531 29055 264537
rect 38565 264537 38577 264540
rect 38611 264537 38623 264571
rect 252186 264568 252192 264580
rect 252147 264540 252192 264568
rect 38565 264531 38623 264537
rect 252186 264528 252192 264540
rect 252244 264528 252250 264580
rect 259178 264568 259184 264580
rect 259139 264540 259184 264568
rect 259178 264528 259184 264540
rect 259236 264528 259242 264580
rect 278041 264571 278099 264577
rect 278041 264537 278053 264571
rect 278087 264568 278099 264571
rect 284662 264568 284668 264580
rect 278087 264540 284668 264568
rect 278087 264537 278099 264540
rect 278041 264531 278099 264537
rect 284662 264528 284668 264540
rect 284720 264528 284726 264580
rect 161106 264460 161112 264512
rect 161164 264500 161170 264512
rect 284478 264500 284484 264512
rect 161164 264472 284484 264500
rect 161164 264460 161170 264472
rect 284478 264460 284484 264472
rect 284536 264460 284542 264512
rect 4985 264435 5043 264441
rect 4985 264401 4997 264435
rect 5031 264432 5043 264435
rect 9677 264435 9735 264441
rect 9677 264432 9689 264435
rect 5031 264404 9689 264432
rect 5031 264401 5043 264404
rect 4985 264395 5043 264401
rect 9677 264401 9689 264404
rect 9723 264401 9735 264435
rect 28997 264435 29055 264441
rect 28997 264432 29009 264435
rect 9677 264395 9735 264401
rect 23308 264404 29009 264432
rect 19245 264367 19303 264373
rect 19245 264333 19257 264367
rect 19291 264364 19303 264367
rect 22005 264367 22063 264373
rect 22005 264364 22017 264367
rect 19291 264336 22017 264364
rect 19291 264333 19303 264336
rect 19245 264327 19303 264333
rect 22005 264333 22017 264336
rect 22051 264333 22063 264367
rect 22005 264327 22063 264333
rect 22097 264367 22155 264373
rect 22097 264333 22109 264367
rect 22143 264364 22155 264367
rect 23308 264364 23336 264404
rect 28997 264401 29009 264404
rect 29043 264401 29055 264435
rect 132862 264432 132868 264444
rect 28997 264395 29055 264401
rect 125520 264404 132868 264432
rect 22143 264336 23336 264364
rect 38565 264367 38623 264373
rect 22143 264333 22155 264336
rect 22097 264327 22155 264333
rect 38565 264333 38577 264367
rect 38611 264364 38623 264367
rect 41417 264367 41475 264373
rect 41417 264364 41429 264367
rect 38611 264336 41429 264364
rect 38611 264333 38623 264336
rect 38565 264327 38623 264333
rect 41417 264333 41429 264336
rect 41463 264333 41475 264367
rect 41417 264327 41475 264333
rect 41509 264367 41567 264373
rect 41509 264333 41521 264367
rect 41555 264364 41567 264367
rect 48317 264367 48375 264373
rect 41555 264336 48268 264364
rect 41555 264333 41567 264336
rect 41509 264327 41567 264333
rect 48240 264296 48268 264336
rect 48317 264333 48329 264367
rect 48363 264333 48375 264367
rect 48317 264327 48375 264333
rect 67637 264367 67695 264373
rect 67637 264333 67649 264367
rect 67683 264364 67695 264367
rect 72421 264367 72479 264373
rect 72421 264364 72433 264367
rect 67683 264336 72433 264364
rect 67683 264333 67695 264336
rect 67637 264327 67695 264333
rect 72421 264333 72433 264336
rect 72467 264333 72479 264367
rect 106277 264367 106335 264373
rect 106277 264364 106289 264367
rect 72421 264327 72479 264333
rect 99576 264336 106289 264364
rect 48332 264296 48360 264327
rect 81434 264296 81440 264308
rect 48240 264268 48360 264296
rect 81395 264268 81440 264296
rect 81434 264256 81440 264268
rect 81492 264256 81498 264308
rect 85574 264296 85580 264308
rect 85535 264268 85580 264296
rect 85574 264256 85580 264268
rect 85632 264256 85638 264308
rect 87414 264296 87420 264308
rect 87375 264268 87420 264296
rect 87414 264256 87420 264268
rect 87472 264256 87478 264308
rect 89717 264299 89775 264305
rect 89717 264265 89729 264299
rect 89763 264296 89775 264299
rect 99285 264299 99343 264305
rect 99285 264296 99297 264299
rect 89763 264268 99297 264296
rect 89763 264265 89775 264268
rect 89717 264259 89775 264265
rect 99285 264265 99297 264268
rect 99331 264265 99343 264299
rect 99285 264259 99343 264265
rect 99377 264299 99435 264305
rect 99377 264265 99389 264299
rect 99423 264296 99435 264299
rect 99576 264296 99604 264336
rect 106277 264333 106289 264336
rect 106323 264333 106335 264367
rect 125520 264364 125548 264404
rect 132862 264392 132868 264404
rect 132920 264392 132926 264444
rect 208394 264392 208400 264444
rect 208452 264432 208458 264444
rect 278041 264435 278099 264441
rect 278041 264432 278053 264435
rect 208452 264404 278053 264432
rect 208452 264392 208458 264404
rect 278041 264401 278053 264404
rect 278087 264401 278099 264435
rect 278041 264395 278099 264401
rect 106277 264327 106335 264333
rect 118528 264336 125548 264364
rect 108666 264296 108672 264308
rect 99423 264268 99604 264296
rect 108627 264268 108672 264296
rect 99423 264265 99435 264268
rect 99377 264259 99435 264265
rect 108666 264256 108672 264268
rect 108724 264256 108730 264308
rect 67637 264231 67695 264237
rect 67637 264228 67649 264231
rect 51092 264200 67649 264228
rect 48317 264163 48375 264169
rect 48317 264129 48329 264163
rect 48363 264160 48375 264163
rect 51092 264160 51120 264200
rect 67637 264197 67649 264200
rect 67683 264197 67695 264231
rect 67637 264191 67695 264197
rect 72421 264231 72479 264237
rect 72421 264197 72433 264231
rect 72467 264228 72479 264231
rect 115845 264231 115903 264237
rect 72467 264200 80100 264228
rect 72467 264197 72479 264200
rect 72421 264191 72479 264197
rect 48363 264132 51120 264160
rect 80072 264160 80100 264200
rect 115845 264197 115857 264231
rect 115891 264228 115903 264231
rect 118528 264228 118556 264336
rect 136450 264324 136456 264376
rect 136508 264364 136514 264376
rect 136508 264336 144500 264364
rect 136508 264324 136514 264336
rect 132310 264256 132316 264308
rect 132368 264256 132374 264308
rect 133506 264296 133512 264308
rect 133467 264268 133512 264296
rect 133506 264256 133512 264268
rect 133564 264256 133570 264308
rect 134426 264296 134432 264308
rect 134387 264268 134432 264296
rect 134426 264256 134432 264268
rect 134484 264256 134490 264308
rect 144362 264256 144368 264308
rect 144420 264256 144426 264308
rect 115891 264200 118556 264228
rect 115891 264197 115903 264200
rect 115845 264191 115903 264197
rect 89717 264163 89775 264169
rect 89717 264160 89729 264163
rect 80072 264132 89729 264160
rect 48363 264129 48375 264132
rect 48317 264123 48375 264129
rect 89717 264129 89729 264132
rect 89763 264129 89775 264163
rect 89717 264123 89775 264129
rect 106277 264095 106335 264101
rect 106277 264061 106289 264095
rect 106323 264092 106335 264095
rect 115845 264095 115903 264101
rect 115845 264092 115857 264095
rect 106323 264064 115857 264092
rect 106323 264061 106335 264064
rect 106277 264055 106335 264061
rect 115845 264061 115857 264064
rect 115891 264061 115903 264095
rect 115845 264055 115903 264061
rect 132328 263956 132356 264256
rect 144380 264024 144408 264256
rect 144472 264160 144500 264336
rect 226242 264324 226248 264376
rect 226300 264364 226306 264376
rect 229741 264367 229799 264373
rect 229741 264364 229753 264367
rect 226300 264336 229753 264364
rect 226300 264324 226306 264336
rect 229741 264333 229753 264336
rect 229787 264333 229799 264367
rect 229741 264327 229799 264333
rect 242250 264324 242256 264376
rect 242308 264364 242314 264376
rect 300854 264364 300860 264376
rect 242308 264336 300860 264364
rect 242308 264324 242314 264336
rect 300854 264324 300860 264336
rect 300912 264324 300918 264376
rect 147674 264296 147680 264308
rect 147635 264268 147680 264296
rect 147674 264256 147680 264268
rect 147732 264256 147738 264308
rect 173802 264296 173808 264308
rect 173763 264268 173808 264296
rect 173802 264256 173808 264268
rect 173860 264256 173866 264308
rect 202690 264296 202696 264308
rect 202651 264268 202696 264296
rect 202690 264256 202696 264268
rect 202748 264256 202754 264308
rect 218514 264256 218520 264308
rect 218572 264256 218578 264308
rect 224402 264296 224408 264308
rect 224363 264268 224408 264296
rect 224402 264256 224408 264268
rect 224460 264256 224466 264308
rect 277949 264299 278007 264305
rect 277949 264296 277961 264299
rect 224512 264268 277961 264296
rect 218532 264228 218560 264256
rect 224512 264228 224540 264268
rect 277949 264265 277961 264268
rect 277995 264265 278007 264299
rect 278682 264296 278688 264308
rect 278643 264268 278688 264296
rect 277949 264259 278007 264265
rect 278682 264256 278688 264268
rect 278740 264256 278746 264308
rect 279786 264256 279792 264308
rect 279844 264296 279850 264308
rect 280798 264296 280804 264308
rect 279844 264268 280804 264296
rect 279844 264256 279850 264268
rect 280798 264256 280804 264268
rect 280856 264256 280862 264308
rect 218532 264200 224540 264228
rect 229741 264231 229799 264237
rect 229741 264197 229753 264231
rect 229787 264228 229799 264231
rect 492674 264228 492680 264240
rect 229787 264200 492680 264228
rect 229787 264197 229799 264200
rect 229741 264191 229799 264197
rect 492674 264188 492680 264200
rect 492732 264188 492738 264240
rect 296714 264160 296720 264172
rect 144472 264132 296720 264160
rect 296714 264120 296720 264132
rect 296772 264120 296778 264172
rect 278685 264095 278743 264101
rect 278685 264061 278697 264095
rect 278731 264092 278743 264095
rect 498194 264092 498200 264104
rect 278731 264064 498200 264092
rect 278731 264061 278743 264064
rect 278685 264055 278743 264061
rect 498194 264052 498200 264064
rect 498252 264052 498258 264104
rect 369854 264024 369860 264036
rect 144380 263996 369860 264024
rect 369854 263984 369860 263996
rect 369912 263984 369918 264036
rect 361574 263956 361580 263968
rect 132328 263928 361580 263956
rect 361574 263916 361580 263928
rect 361632 263916 361638 263968
rect 133509 263891 133567 263897
rect 133509 263857 133521 263891
rect 133555 263888 133567 263891
rect 375374 263888 375380 263900
rect 133555 263860 375380 263888
rect 133555 263857 133567 263860
rect 133509 263851 133567 263857
rect 375374 263848 375380 263860
rect 375432 263848 375438 263900
rect 56502 263780 56508 263832
rect 56560 263820 56566 263832
rect 81437 263823 81495 263829
rect 81437 263820 81449 263823
rect 56560 263792 81449 263820
rect 56560 263780 56566 263792
rect 81437 263789 81449 263792
rect 81483 263789 81495 263823
rect 81437 263783 81495 263789
rect 202693 263823 202751 263829
rect 202693 263789 202705 263823
rect 202739 263820 202751 263823
rect 451274 263820 451280 263832
rect 202739 263792 451280 263820
rect 202739 263789 202751 263792
rect 202693 263783 202751 263789
rect 451274 263780 451280 263792
rect 451332 263780 451338 263832
rect 56410 263712 56416 263764
rect 56468 263752 56474 263764
rect 85577 263755 85635 263761
rect 85577 263752 85589 263755
rect 56468 263724 85589 263752
rect 56468 263712 56474 263724
rect 85577 263721 85589 263724
rect 85623 263721 85635 263755
rect 85577 263715 85635 263721
rect 134429 263755 134487 263761
rect 134429 263721 134441 263755
rect 134475 263752 134487 263755
rect 390554 263752 390560 263764
rect 134475 263724 390560 263752
rect 134475 263721 134487 263724
rect 134429 263715 134487 263721
rect 390554 263712 390560 263724
rect 390612 263712 390618 263764
rect 55030 263644 55036 263696
rect 55088 263684 55094 263696
rect 87417 263687 87475 263693
rect 87417 263684 87429 263687
rect 55088 263656 87429 263684
rect 55088 263644 55094 263656
rect 87417 263653 87429 263656
rect 87463 263653 87475 263687
rect 87417 263647 87475 263653
rect 108669 263687 108727 263693
rect 108669 263653 108681 263687
rect 108715 263684 108727 263687
rect 368474 263684 368480 263696
rect 108715 263656 368480 263684
rect 108715 263653 108727 263656
rect 108669 263647 108727 263653
rect 368474 263644 368480 263656
rect 368532 263644 368538 263696
rect 53650 263576 53656 263628
rect 53708 263616 53714 263628
rect 147677 263619 147735 263625
rect 147677 263616 147689 263619
rect 53708 263588 147689 263616
rect 53708 263576 53714 263588
rect 147677 263585 147689 263588
rect 147723 263585 147735 263619
rect 147677 263579 147735 263585
rect 259181 263619 259239 263625
rect 259181 263585 259193 263619
rect 259227 263616 259239 263619
rect 527174 263616 527180 263628
rect 259227 263588 527180 263616
rect 259227 263585 259239 263588
rect 259181 263579 259239 263585
rect 527174 263576 527180 263588
rect 527232 263576 527238 263628
rect 281350 263508 281356 263560
rect 281408 263548 281414 263560
rect 288434 263548 288440 263560
rect 281408 263520 288440 263548
rect 281408 263508 281414 263520
rect 288434 263508 288440 263520
rect 288492 263508 288498 263560
rect 429378 263548 429384 263560
rect 429339 263520 429384 263548
rect 429378 263508 429384 263520
rect 429436 263508 429442 263560
rect 282178 263440 282184 263492
rect 282236 263480 282242 263492
rect 282454 263480 282460 263492
rect 282236 263452 282460 263480
rect 282236 263440 282242 263452
rect 282454 263440 282460 263452
rect 282512 263440 282518 263492
rect 280982 263168 280988 263220
rect 281040 263208 281046 263220
rect 556154 263208 556160 263220
rect 281040 263180 556160 263208
rect 281040 263168 281046 263180
rect 556154 263168 556160 263180
rect 556212 263168 556218 263220
rect 271785 263143 271843 263149
rect 271785 263109 271797 263143
rect 271831 263140 271843 263143
rect 499574 263140 499580 263152
rect 271831 263112 499580 263140
rect 271831 263109 271843 263112
rect 271785 263103 271843 263109
rect 499574 263100 499580 263112
rect 499632 263100 499638 263152
rect 252189 263075 252247 263081
rect 252189 263041 252201 263075
rect 252235 263072 252247 263075
rect 285858 263072 285864 263084
rect 252235 263044 285864 263072
rect 252235 263041 252247 263044
rect 252189 263035 252247 263041
rect 285858 263032 285864 263044
rect 285916 263032 285922 263084
rect 173805 263007 173863 263013
rect 173805 262973 173817 263007
rect 173851 263004 173863 263007
rect 281074 263004 281080 263016
rect 173851 262976 281080 263004
rect 173851 262973 173863 262976
rect 173805 262967 173863 262973
rect 281074 262964 281080 262976
rect 281132 262964 281138 263016
rect 224405 262939 224463 262945
rect 224405 262905 224417 262939
rect 224451 262936 224463 262939
rect 357434 262936 357440 262948
rect 224451 262908 357440 262936
rect 224451 262905 224463 262908
rect 224405 262899 224463 262905
rect 357434 262896 357440 262908
rect 357492 262896 357498 262948
rect 263597 262871 263655 262877
rect 263597 262837 263609 262871
rect 263643 262868 263655 262871
rect 445754 262868 445760 262880
rect 263643 262840 445760 262868
rect 263643 262837 263655 262840
rect 263597 262831 263655 262837
rect 445754 262828 445760 262840
rect 445812 262828 445818 262880
rect 60274 262760 60280 262812
rect 60332 262800 60338 262812
rect 286594 262800 286600 262812
rect 60332 262772 286600 262800
rect 60332 262760 60338 262772
rect 286594 262760 286600 262772
rect 286652 262760 286658 262812
rect 282362 261604 282368 261656
rect 282420 261644 282426 261656
rect 296806 261644 296812 261656
rect 282420 261616 296812 261644
rect 282420 261604 282426 261616
rect 296806 261604 296812 261616
rect 296864 261604 296870 261656
rect 281166 261536 281172 261588
rect 281224 261576 281230 261588
rect 451366 261576 451372 261588
rect 281224 261548 451372 261576
rect 281224 261536 281230 261548
rect 451366 261536 451372 261548
rect 451424 261536 451430 261588
rect 280982 261468 280988 261520
rect 281040 261508 281046 261520
rect 459554 261508 459560 261520
rect 281040 261480 459560 261508
rect 281040 261468 281046 261480
rect 459554 261468 459560 261480
rect 459612 261468 459618 261520
rect 1302 261400 1308 261452
rect 1360 261440 1366 261452
rect 4985 261443 5043 261449
rect 4985 261440 4997 261443
rect 1360 261412 4997 261440
rect 1360 261400 1366 261412
rect 4985 261409 4997 261412
rect 5031 261409 5043 261443
rect 4985 261403 5043 261409
rect 283190 260856 283196 260908
rect 283248 260896 283254 260908
rect 304258 260896 304264 260908
rect 283248 260868 304264 260896
rect 283248 260856 283254 260868
rect 304258 260856 304264 260868
rect 304316 260856 304322 260908
rect 6178 260788 6184 260840
rect 6236 260828 6242 260840
rect 59354 260828 59360 260840
rect 6236 260800 59360 260828
rect 6236 260788 6242 260800
rect 59354 260788 59360 260800
rect 59412 260788 59418 260840
rect 299474 260788 299480 260840
rect 299532 260828 299538 260840
rect 299658 260828 299664 260840
rect 299532 260800 299664 260828
rect 299532 260788 299538 260800
rect 299658 260788 299664 260800
rect 299716 260788 299722 260840
rect 429378 260788 429384 260840
rect 429436 260828 429442 260840
rect 429565 260831 429623 260837
rect 429565 260828 429577 260831
rect 429436 260800 429577 260828
rect 429436 260788 429442 260800
rect 429565 260797 429577 260800
rect 429611 260797 429623 260831
rect 429565 260791 429623 260797
rect 280890 260176 280896 260228
rect 280948 260216 280954 260228
rect 455414 260216 455420 260228
rect 280948 260188 455420 260216
rect 280948 260176 280954 260188
rect 455414 260176 455420 260188
rect 455472 260176 455478 260228
rect 281258 260108 281264 260160
rect 281316 260148 281322 260160
rect 485774 260148 485780 260160
rect 281316 260120 485780 260148
rect 281316 260108 281322 260120
rect 485774 260108 485780 260120
rect 485832 260108 485838 260160
rect 283098 258748 283104 258800
rect 283156 258788 283162 258800
rect 306374 258788 306380 258800
rect 283156 258760 306380 258788
rect 283156 258748 283162 258760
rect 306374 258748 306380 258760
rect 306432 258748 306438 258800
rect 281994 258680 282000 258732
rect 282052 258720 282058 258732
rect 367094 258720 367100 258732
rect 282052 258692 367100 258720
rect 282052 258680 282058 258692
rect 367094 258680 367100 258692
rect 367152 258680 367158 258732
rect 282270 257320 282276 257372
rect 282328 257360 282334 257372
rect 467834 257360 467840 257372
rect 282328 257332 467840 257360
rect 282328 257320 282334 257332
rect 467834 257320 467840 257332
rect 467892 257320 467898 257372
rect 283558 255960 283564 256012
rect 283616 256000 283622 256012
rect 402974 256000 402980 256012
rect 283616 255972 402980 256000
rect 283616 255960 283622 255972
rect 402974 255960 402980 255972
rect 403032 255960 403038 256012
rect 429562 253960 429568 253972
rect 429523 253932 429568 253960
rect 429562 253920 429568 253932
rect 429620 253920 429626 253972
rect 280798 253172 280804 253224
rect 280856 253212 280862 253224
rect 578234 253212 578240 253224
rect 280856 253184 578240 253212
rect 280856 253172 280862 253184
rect 578234 253172 578240 253184
rect 578292 253172 578298 253224
rect 286594 252492 286600 252544
rect 286652 252532 286658 252544
rect 579798 252532 579804 252544
rect 286652 252504 579804 252532
rect 286652 252492 286658 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 4062 251200 4068 251252
rect 4120 251240 4126 251252
rect 8938 251240 8944 251252
rect 4120 251212 8944 251240
rect 4120 251200 4126 251212
rect 8938 251200 8944 251212
rect 8996 251200 9002 251252
rect 284110 251200 284116 251252
rect 284168 251240 284174 251252
rect 332594 251240 332600 251252
rect 284168 251212 332600 251240
rect 284168 251200 284174 251212
rect 332594 251200 332600 251212
rect 332652 251200 332658 251252
rect 284202 251132 284208 251184
rect 284260 251172 284266 251184
rect 304350 251172 304356 251184
rect 284260 251144 304356 251172
rect 284260 251132 284266 251144
rect 304350 251132 304356 251144
rect 304408 251132 304414 251184
rect 284202 248412 284208 248464
rect 284260 248452 284266 248464
rect 302234 248452 302240 248464
rect 284260 248424 302240 248452
rect 284260 248412 284266 248424
rect 302234 248412 302240 248424
rect 302292 248412 302298 248464
rect 284202 245624 284208 245676
rect 284260 245664 284266 245676
rect 311894 245664 311900 245676
rect 284260 245636 311900 245664
rect 284260 245624 284266 245636
rect 311894 245624 311900 245636
rect 311952 245624 311958 245676
rect 284202 244264 284208 244316
rect 284260 244304 284266 244316
rect 535454 244304 535460 244316
rect 284260 244276 535460 244304
rect 284260 244264 284266 244276
rect 535454 244264 535460 244276
rect 535512 244264 535518 244316
rect 542354 244196 542360 244248
rect 542412 244236 542418 244248
rect 542630 244236 542636 244248
rect 542412 244208 542636 244236
rect 542412 244196 542418 244208
rect 542630 244196 542636 244208
rect 542688 244196 542694 244248
rect 287974 243516 287980 243568
rect 288032 243556 288038 243568
rect 400214 243556 400220 243568
rect 288032 243528 400220 243556
rect 288032 243516 288038 243528
rect 400214 243516 400220 243528
rect 400272 243516 400278 243568
rect 283834 238688 283840 238740
rect 283892 238728 283898 238740
rect 319438 238728 319444 238740
rect 283892 238700 319444 238728
rect 283892 238688 283898 238700
rect 319438 238688 319444 238700
rect 319496 238688 319502 238740
rect 282178 238008 282184 238060
rect 282236 238048 282242 238060
rect 396074 238048 396080 238060
rect 282236 238020 396080 238048
rect 282236 238008 282242 238020
rect 396074 238008 396080 238020
rect 396132 238008 396138 238060
rect 4062 237328 4068 237380
rect 4120 237368 4126 237380
rect 17218 237368 17224 237380
rect 4120 237340 17224 237368
rect 4120 237328 4126 237340
rect 17218 237328 17224 237340
rect 17276 237328 17282 237380
rect 429286 234676 429292 234728
rect 429344 234676 429350 234728
rect 429304 234592 429332 234676
rect 429286 234540 429292 234592
rect 429344 234540 429350 234592
rect 284202 233248 284208 233300
rect 284260 233288 284266 233300
rect 308398 233288 308404 233300
rect 284260 233260 308404 233288
rect 284260 233248 284266 233260
rect 308398 233248 308404 233260
rect 308456 233248 308462 233300
rect 7926 231820 7932 231872
rect 7984 231860 7990 231872
rect 8018 231860 8024 231872
rect 7984 231832 8024 231860
rect 7984 231820 7990 231832
rect 8018 231820 8024 231832
rect 8076 231820 8082 231872
rect 299474 231820 299480 231872
rect 299532 231860 299538 231872
rect 299750 231860 299756 231872
rect 299532 231832 299756 231860
rect 299532 231820 299538 231832
rect 299750 231820 299756 231832
rect 299808 231820 299814 231872
rect 542538 231820 542544 231872
rect 542596 231860 542602 231872
rect 542722 231860 542728 231872
rect 542596 231832 542728 231860
rect 542596 231820 542602 231832
rect 542722 231820 542728 231832
rect 542780 231820 542786 231872
rect 429286 231792 429292 231804
rect 429247 231764 429292 231792
rect 429286 231752 429292 231764
rect 429344 231752 429350 231804
rect 284110 228556 284116 228608
rect 284168 228596 284174 228608
rect 286502 228596 286508 228608
rect 284168 228568 286508 228596
rect 284168 228556 284174 228568
rect 286502 228556 286508 228568
rect 286560 228556 286566 228608
rect 284202 226312 284208 226364
rect 284260 226352 284266 226364
rect 467098 226352 467104 226364
rect 284260 226324 467104 226352
rect 284260 226312 284266 226324
rect 467098 226312 467104 226324
rect 467156 226312 467162 226364
rect 284202 224952 284208 225004
rect 284260 224992 284266 225004
rect 497458 224992 497464 225004
rect 284260 224964 497464 224992
rect 284260 224952 284266 224964
rect 497458 224952 497464 224964
rect 497516 224952 497522 225004
rect 3602 223524 3608 223576
rect 3660 223564 3666 223576
rect 59354 223564 59360 223576
rect 3660 223536 59360 223564
rect 3660 223524 3666 223536
rect 59354 223524 59360 223536
rect 59412 223524 59418 223576
rect 2958 223456 2964 223508
rect 3016 223496 3022 223508
rect 19978 223496 19984 223508
rect 3016 223468 19984 223496
rect 3016 223456 3022 223468
rect 19978 223456 19984 223468
rect 20036 223456 20042 223508
rect 429289 222207 429347 222213
rect 429289 222173 429301 222207
rect 429335 222204 429347 222207
rect 429470 222204 429476 222216
rect 429335 222176 429476 222204
rect 429335 222173 429347 222176
rect 429289 222167 429347 222173
rect 429470 222164 429476 222176
rect 429528 222164 429534 222216
rect 542354 222164 542360 222216
rect 542412 222204 542418 222216
rect 542630 222204 542636 222216
rect 542412 222176 542636 222204
rect 542412 222164 542418 222176
rect 542630 222164 542636 222176
rect 542688 222164 542694 222216
rect 8018 222136 8024 222148
rect 7979 222108 8024 222136
rect 8018 222096 8024 222108
rect 8076 222096 8082 222148
rect 53558 220804 53564 220856
rect 53616 220844 53622 220856
rect 59354 220844 59360 220856
rect 53616 220816 59360 220844
rect 53616 220804 53622 220816
rect 59354 220804 59360 220816
rect 59412 220804 59418 220856
rect 53466 216656 53472 216708
rect 53524 216696 53530 216708
rect 59446 216696 59452 216708
rect 53524 216668 59452 216696
rect 53524 216656 53530 216668
rect 59446 216656 59452 216668
rect 59504 216656 59510 216708
rect 284202 216656 284208 216708
rect 284260 216696 284266 216708
rect 385678 216696 385684 216708
rect 284260 216668 385684 216696
rect 284260 216656 284266 216668
rect 385678 216656 385684 216668
rect 385736 216656 385742 216708
rect 14550 216588 14556 216640
rect 14608 216628 14614 216640
rect 59354 216628 59360 216640
rect 14608 216600 59360 216628
rect 14608 216588 14614 216600
rect 59354 216588 59360 216600
rect 59412 216588 59418 216640
rect 284202 215296 284208 215348
rect 284260 215336 284266 215348
rect 514018 215336 514024 215348
rect 284260 215308 514024 215336
rect 284260 215296 284266 215308
rect 514018 215296 514024 215308
rect 514076 215296 514082 215348
rect 8021 215203 8079 215209
rect 8021 215169 8033 215203
rect 8067 215200 8079 215203
rect 8110 215200 8116 215212
rect 8067 215172 8116 215200
rect 8067 215169 8079 215172
rect 8021 215163 8079 215169
rect 8110 215160 8116 215172
rect 8168 215160 8174 215212
rect 429286 215160 429292 215212
rect 429344 215200 429350 215212
rect 429470 215200 429476 215212
rect 429344 215172 429476 215200
rect 429344 215160 429350 215172
rect 429470 215160 429476 215172
rect 429528 215160 429534 215212
rect 54938 213936 54944 213988
rect 54996 213976 55002 213988
rect 59354 213976 59360 213988
rect 54996 213948 59360 213976
rect 54996 213936 55002 213948
rect 59354 213936 59360 213948
rect 59412 213936 59418 213988
rect 299474 212576 299480 212628
rect 299532 212616 299538 212628
rect 299750 212616 299756 212628
rect 299532 212588 299756 212616
rect 299532 212576 299538 212588
rect 299750 212576 299756 212588
rect 299808 212576 299814 212628
rect 56134 212508 56140 212560
rect 56192 212548 56198 212560
rect 59354 212548 59360 212560
rect 56192 212520 59360 212548
rect 56192 212508 56198 212520
rect 59354 212508 59360 212520
rect 59412 212508 59418 212560
rect 284202 212508 284208 212560
rect 284260 212548 284266 212560
rect 331214 212548 331220 212560
rect 284260 212520 331220 212548
rect 284260 212508 284266 212520
rect 331214 212508 331220 212520
rect 331272 212508 331278 212560
rect 284202 211148 284208 211200
rect 284260 211188 284266 211200
rect 462314 211188 462320 211200
rect 284260 211160 462320 211188
rect 284260 211148 284266 211160
rect 462314 211148 462320 211160
rect 462372 211148 462378 211200
rect 280890 209788 280896 209840
rect 280948 209828 280954 209840
rect 281166 209828 281172 209840
rect 280948 209800 281172 209828
rect 280948 209788 280954 209800
rect 281166 209788 281172 209800
rect 281224 209788 281230 209840
rect 280798 209760 280804 209772
rect 280759 209732 280804 209760
rect 280798 209720 280804 209732
rect 280856 209720 280862 209772
rect 284110 207000 284116 207052
rect 284168 207040 284174 207052
rect 478874 207040 478880 207052
rect 284168 207012 478880 207040
rect 284168 207000 284174 207012
rect 478874 207000 478880 207012
rect 478932 207000 478938 207052
rect 8110 205748 8116 205760
rect 7944 205720 8116 205748
rect 7944 205624 7972 205720
rect 8110 205708 8116 205720
rect 8168 205708 8174 205760
rect 53374 205640 53380 205692
rect 53432 205680 53438 205692
rect 59354 205680 59360 205692
rect 53432 205652 59360 205680
rect 53432 205640 53438 205652
rect 59354 205640 59360 205652
rect 59412 205640 59418 205692
rect 7926 205572 7932 205624
rect 7984 205572 7990 205624
rect 429286 205572 429292 205624
rect 429344 205612 429350 205624
rect 429470 205612 429476 205624
rect 429344 205584 429476 205612
rect 429344 205572 429350 205584
rect 429470 205572 429476 205584
rect 429528 205572 429534 205624
rect 284202 204348 284208 204400
rect 284260 204388 284266 204400
rect 305638 204388 305644 204400
rect 284260 204360 305644 204388
rect 284260 204348 284266 204360
rect 305638 204348 305644 204360
rect 305696 204348 305702 204400
rect 304350 204280 304356 204332
rect 304408 204320 304414 204332
rect 579890 204320 579896 204332
rect 304408 204292 579896 204320
rect 304408 204280 304414 204292
rect 579890 204280 579896 204292
rect 579948 204280 579954 204332
rect 54846 202852 54852 202904
rect 54904 202892 54910 202904
rect 59354 202892 59360 202904
rect 54904 202864 59360 202892
rect 54904 202852 54910 202864
rect 59354 202852 59360 202864
rect 59412 202852 59418 202904
rect 542538 202852 542544 202904
rect 542596 202892 542602 202904
rect 542630 202892 542636 202904
rect 542596 202864 542636 202892
rect 542596 202852 542602 202864
rect 542630 202852 542636 202864
rect 542688 202852 542694 202904
rect 299658 202824 299664 202836
rect 299619 202796 299664 202824
rect 299658 202784 299664 202796
rect 299716 202784 299722 202836
rect 429470 202824 429476 202836
rect 429431 202796 429476 202824
rect 429470 202784 429476 202796
rect 429528 202784 429534 202836
rect 284202 201492 284208 201544
rect 284260 201532 284266 201544
rect 337378 201532 337384 201544
rect 284260 201504 337384 201532
rect 284260 201492 284266 201504
rect 337378 201492 337384 201504
rect 337436 201492 337442 201544
rect 7926 201464 7932 201476
rect 7887 201436 7932 201464
rect 7926 201424 7932 201436
rect 7984 201424 7990 201476
rect 280801 200175 280859 200181
rect 280801 200141 280813 200175
rect 280847 200172 280859 200175
rect 280982 200172 280988 200184
rect 280847 200144 280988 200172
rect 280847 200141 280859 200144
rect 280801 200135 280859 200141
rect 280982 200132 280988 200144
rect 281040 200132 281046 200184
rect 24118 200064 24124 200116
rect 24176 200104 24182 200116
rect 59354 200104 59360 200116
rect 24176 200076 59360 200104
rect 24176 200064 24182 200076
rect 59354 200064 59360 200076
rect 59412 200064 59418 200116
rect 280982 200036 280988 200048
rect 280943 200008 280988 200036
rect 280982 199996 280988 200008
rect 281040 199996 281046 200048
rect 284202 198704 284208 198756
rect 284260 198744 284266 198756
rect 430574 198744 430580 198756
rect 284260 198716 430580 198744
rect 284260 198704 284266 198716
rect 430574 198704 430580 198716
rect 430632 198704 430638 198756
rect 542630 195984 542636 196036
rect 542688 195984 542694 196036
rect 542648 195956 542676 195984
rect 542722 195956 542728 195968
rect 542648 195928 542728 195956
rect 542722 195916 542728 195928
rect 542780 195916 542786 195968
rect 27614 194488 27620 194540
rect 27672 194528 27678 194540
rect 37182 194528 37188 194540
rect 27672 194500 37188 194528
rect 27672 194488 27678 194500
rect 37182 194488 37188 194500
rect 37240 194488 37246 194540
rect 299661 193307 299719 193313
rect 299661 193273 299673 193307
rect 299707 193304 299719 193307
rect 299750 193304 299756 193316
rect 299707 193276 299756 193304
rect 299707 193273 299719 193276
rect 299661 193267 299719 193273
rect 299750 193264 299756 193276
rect 299808 193264 299814 193316
rect 429473 193307 429531 193313
rect 429473 193273 429485 193307
rect 429519 193304 429531 193307
rect 429562 193304 429568 193316
rect 429519 193276 429568 193304
rect 429519 193273 429531 193276
rect 429473 193267 429531 193273
rect 429562 193264 429568 193276
rect 429620 193264 429626 193316
rect 53282 193196 53288 193248
rect 53340 193236 53346 193248
rect 59354 193236 59360 193248
rect 53340 193208 59360 193236
rect 53340 193196 53346 193208
rect 59354 193196 59360 193208
rect 59412 193196 59418 193248
rect 284202 193196 284208 193248
rect 284260 193236 284266 193248
rect 517514 193236 517520 193248
rect 284260 193208 517520 193236
rect 284260 193196 284266 193208
rect 517514 193196 517520 193208
rect 517572 193196 517578 193248
rect 7926 193168 7932 193180
rect 7887 193140 7932 193168
rect 7926 193128 7932 193140
rect 7984 193128 7990 193180
rect 280982 190856 280988 190868
rect 280943 190828 280988 190856
rect 280982 190816 280988 190828
rect 281040 190816 281046 190868
rect 3694 188980 3700 189032
rect 3752 189020 3758 189032
rect 59354 189020 59360 189032
rect 3752 188992 59360 189020
rect 3752 188980 3758 188992
rect 59354 188980 59360 188992
rect 59412 188980 59418 189032
rect 284202 187688 284208 187740
rect 284260 187728 284266 187740
rect 364978 187728 364984 187740
rect 284260 187700 364984 187728
rect 284260 187688 284266 187700
rect 364978 187688 364984 187700
rect 365036 187688 365042 187740
rect 8018 186328 8024 186380
rect 8076 186368 8082 186380
rect 8076 186340 8156 186368
rect 8076 186328 8082 186340
rect 8128 186244 8156 186340
rect 8110 186192 8116 186244
rect 8168 186192 8174 186244
rect 542538 183540 542544 183592
rect 542596 183580 542602 183592
rect 542814 183580 542820 183592
rect 542596 183552 542820 183580
rect 542596 183540 542602 183552
rect 542814 183540 542820 183552
rect 542872 183540 542878 183592
rect 429470 183512 429476 183524
rect 429431 183484 429476 183512
rect 429470 183472 429476 183484
rect 429528 183472 429534 183524
rect 57606 182180 57612 182232
rect 57664 182220 57670 182232
rect 59906 182220 59912 182232
rect 57664 182192 59912 182220
rect 57664 182180 57670 182192
rect 59906 182180 59912 182192
rect 59964 182180 59970 182232
rect 284202 182180 284208 182232
rect 284260 182220 284266 182232
rect 292574 182220 292580 182232
rect 284260 182192 292580 182220
rect 284260 182180 284266 182192
rect 292574 182180 292580 182192
rect 292632 182180 292638 182232
rect 293310 182112 293316 182164
rect 293368 182152 293374 182164
rect 580166 182152 580172 182164
rect 293368 182124 580172 182152
rect 293368 182112 293374 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 53190 180820 53196 180872
rect 53248 180860 53254 180872
rect 59354 180860 59360 180872
rect 53248 180832 59360 180860
rect 53248 180820 53254 180832
rect 59354 180820 59360 180832
rect 59412 180820 59418 180872
rect 280982 179324 280988 179376
rect 281040 179364 281046 179376
rect 281442 179364 281448 179376
rect 281040 179336 281448 179364
rect 281040 179324 281046 179336
rect 281442 179324 281448 179336
rect 281500 179324 281506 179376
rect 8110 176740 8116 176792
rect 8168 176740 8174 176792
rect 8018 176536 8024 176588
rect 8076 176576 8082 176588
rect 8128 176576 8156 176740
rect 284202 176672 284208 176724
rect 284260 176712 284266 176724
rect 502978 176712 502984 176724
rect 284260 176684 502984 176712
rect 284260 176672 284266 176684
rect 502978 176672 502984 176684
rect 503036 176672 503042 176724
rect 8076 176548 8156 176576
rect 8076 176536 8082 176548
rect 57514 175244 57520 175296
rect 57572 175284 57578 175296
rect 59538 175284 59544 175296
rect 57572 175256 59544 175284
rect 57572 175244 57578 175256
rect 59538 175244 59544 175256
rect 59596 175244 59602 175296
rect 299474 173952 299480 174004
rect 299532 173992 299538 174004
rect 299750 173992 299756 174004
rect 299532 173964 299756 173992
rect 299532 173952 299538 173964
rect 299750 173952 299756 173964
rect 299808 173952 299814 174004
rect 429473 173995 429531 174001
rect 429473 173961 429485 173995
rect 429519 173992 429531 173995
rect 429562 173992 429568 174004
rect 429519 173964 429568 173992
rect 429519 173961 429531 173964
rect 429473 173955 429531 173961
rect 429562 173952 429568 173964
rect 429620 173952 429626 174004
rect 284202 173884 284208 173936
rect 284260 173924 284266 173936
rect 477494 173924 477500 173936
rect 284260 173896 477500 173924
rect 284260 173884 284266 173896
rect 477494 173884 477500 173896
rect 477552 173884 477558 173936
rect 542630 173884 542636 173936
rect 542688 173924 542694 173936
rect 542814 173924 542820 173936
rect 542688 173896 542820 173924
rect 542688 173884 542694 173896
rect 542814 173884 542820 173896
rect 542872 173884 542878 173936
rect 280798 171912 280804 171964
rect 280856 171952 280862 171964
rect 281166 171952 281172 171964
rect 280856 171924 281172 171952
rect 280856 171912 280862 171924
rect 281166 171912 281172 171924
rect 281224 171912 281230 171964
rect 284202 171096 284208 171148
rect 284260 171136 284266 171148
rect 447134 171136 447140 171148
rect 284260 171108 447140 171136
rect 284260 171096 284266 171108
rect 447134 171096 447140 171108
rect 447192 171096 447198 171148
rect 285306 169736 285312 169788
rect 285364 169776 285370 169788
rect 580166 169776 580172 169788
rect 285364 169748 580172 169776
rect 285364 169736 285370 169748
rect 580166 169736 580172 169748
rect 580224 169736 580230 169788
rect 542354 169056 542360 169108
rect 542412 169096 542418 169108
rect 542630 169096 542636 169108
rect 542412 169068 542636 169096
rect 542412 169056 542418 169068
rect 542630 169056 542636 169068
rect 542688 169056 542694 169108
rect 15838 168308 15844 168360
rect 15896 168348 15902 168360
rect 59354 168348 59360 168360
rect 15896 168320 59360 168348
rect 15896 168308 15902 168320
rect 59354 168308 59360 168320
rect 59412 168308 59418 168360
rect 281258 166880 281264 166932
rect 281316 166920 281322 166932
rect 281442 166920 281448 166932
rect 281316 166892 281448 166920
rect 281316 166880 281322 166892
rect 281442 166880 281448 166892
rect 281500 166880 281506 166932
rect 3326 165520 3332 165572
rect 3384 165560 3390 165572
rect 6270 165560 6276 165572
rect 3384 165532 6276 165560
rect 3384 165520 3390 165532
rect 6270 165520 6276 165532
rect 6328 165520 6334 165572
rect 13078 165520 13084 165572
rect 13136 165560 13142 165572
rect 59354 165560 59360 165572
rect 13136 165532 59360 165560
rect 13136 165520 13142 165532
rect 59354 165520 59360 165532
rect 59412 165520 59418 165572
rect 283834 164228 283840 164280
rect 283892 164268 283898 164280
rect 501598 164268 501604 164280
rect 283892 164240 501604 164268
rect 283892 164228 283898 164240
rect 501598 164228 501604 164240
rect 501656 164228 501662 164280
rect 8018 164160 8024 164212
rect 8076 164200 8082 164212
rect 8110 164200 8116 164212
rect 8076 164172 8116 164200
rect 8076 164160 8082 164172
rect 8110 164160 8116 164172
rect 8168 164160 8174 164212
rect 299474 164160 299480 164212
rect 299532 164200 299538 164212
rect 299658 164200 299664 164212
rect 299532 164172 299664 164200
rect 299532 164160 299538 164172
rect 299658 164160 299664 164172
rect 299716 164160 299722 164212
rect 429378 164200 429384 164212
rect 429339 164172 429384 164200
rect 429378 164160 429384 164172
rect 429436 164160 429442 164212
rect 283834 162868 283840 162920
rect 283892 162908 283898 162920
rect 371878 162908 371884 162920
rect 283892 162880 371884 162908
rect 283892 162868 283898 162880
rect 371878 162868 371884 162880
rect 371936 162868 371942 162920
rect 280798 162120 280804 162172
rect 280856 162160 280862 162172
rect 281258 162160 281264 162172
rect 280856 162132 281264 162160
rect 280856 162120 280862 162132
rect 281258 162120 281264 162132
rect 281316 162120 281322 162172
rect 542354 161372 542360 161424
rect 542412 161412 542418 161424
rect 542630 161412 542636 161424
rect 542412 161384 542636 161412
rect 542412 161372 542418 161384
rect 542630 161372 542636 161384
rect 542688 161372 542694 161424
rect 283374 160080 283380 160132
rect 283432 160120 283438 160132
rect 316034 160120 316040 160132
rect 283432 160092 316040 160120
rect 283432 160080 283438 160092
rect 316034 160080 316040 160092
rect 316092 160080 316098 160132
rect 422938 157360 422944 157412
rect 422996 157400 423002 157412
rect 579890 157400 579896 157412
rect 422996 157372 579896 157400
rect 422996 157360 423002 157372
rect 579890 157360 579896 157372
rect 579948 157360 579954 157412
rect 429378 157332 429384 157344
rect 429339 157304 429384 157332
rect 429378 157292 429384 157304
rect 429436 157292 429442 157344
rect 284018 153212 284024 153264
rect 284076 153252 284082 153264
rect 322290 153252 322296 153264
rect 284076 153224 322296 153252
rect 284076 153212 284082 153224
rect 322290 153212 322296 153224
rect 322348 153212 322354 153264
rect 280798 152600 280804 152652
rect 280856 152640 280862 152652
rect 281166 152640 281172 152652
rect 280856 152612 281172 152640
rect 280856 152600 280862 152612
rect 281166 152600 281172 152612
rect 281224 152600 281230 152652
rect 280798 152396 280804 152448
rect 280856 152436 280862 152448
rect 281258 152436 281264 152448
rect 280856 152408 281264 152436
rect 280856 152396 280862 152408
rect 281258 152396 281264 152408
rect 281316 152396 281322 152448
rect 542354 151784 542360 151836
rect 542412 151824 542418 151836
rect 542630 151824 542636 151836
rect 542412 151796 542636 151824
rect 542412 151784 542418 151796
rect 542630 151784 542636 151796
rect 542688 151784 542694 151836
rect 6178 150424 6184 150476
rect 6236 150464 6242 150476
rect 59354 150464 59360 150476
rect 6236 150436 59360 150464
rect 6236 150424 6242 150436
rect 59354 150424 59360 150436
rect 59412 150424 59418 150476
rect 283834 150356 283840 150408
rect 283892 150396 283898 150408
rect 315298 150396 315304 150408
rect 283892 150368 315304 150396
rect 283892 150356 283898 150368
rect 315298 150356 315304 150368
rect 315356 150356 315362 150408
rect 429286 147636 429292 147688
rect 429344 147676 429350 147688
rect 429470 147676 429476 147688
rect 429344 147648 429476 147676
rect 429344 147636 429350 147648
rect 429470 147636 429476 147648
rect 429528 147636 429534 147688
rect 8018 144848 8024 144900
rect 8076 144888 8082 144900
rect 8110 144888 8116 144900
rect 8076 144860 8116 144888
rect 8076 144848 8082 144860
rect 8110 144848 8116 144860
rect 8168 144848 8174 144900
rect 283834 144848 283840 144900
rect 283892 144888 283898 144900
rect 422938 144888 422944 144900
rect 283892 144860 422944 144888
rect 283892 144848 283898 144860
rect 422938 144848 422944 144860
rect 422996 144848 423002 144900
rect 429378 144888 429384 144900
rect 429339 144860 429384 144888
rect 429378 144848 429384 144860
rect 429436 144848 429442 144900
rect 57422 142604 57428 142656
rect 57480 142644 57486 142656
rect 59354 142644 59360 142656
rect 57480 142616 59360 142644
rect 57480 142604 57486 142616
rect 59354 142604 59360 142616
rect 59412 142604 59418 142656
rect 283834 142128 283840 142180
rect 283892 142168 283898 142180
rect 372614 142168 372620 142180
rect 283892 142140 372620 142168
rect 283892 142128 283898 142140
rect 372614 142128 372620 142140
rect 372672 142128 372678 142180
rect 284202 142060 284208 142112
rect 284260 142100 284266 142112
rect 313918 142100 313924 142112
rect 284260 142072 313924 142100
rect 284260 142060 284266 142072
rect 313918 142060 313924 142072
rect 313976 142060 313982 142112
rect 542354 142060 542360 142112
rect 542412 142100 542418 142112
rect 542630 142100 542636 142112
rect 542412 142072 542636 142100
rect 542412 142060 542418 142072
rect 542630 142060 542636 142072
rect 542688 142060 542694 142112
rect 429378 137952 429384 137964
rect 429339 137924 429384 137952
rect 429378 137912 429384 137924
rect 429436 137912 429442 137964
rect 283742 136620 283748 136672
rect 283800 136660 283806 136672
rect 426434 136660 426440 136672
rect 283800 136632 426440 136660
rect 283800 136620 283806 136632
rect 426434 136620 426440 136632
rect 426492 136620 426498 136672
rect 3970 135260 3976 135312
rect 4028 135300 4034 135312
rect 53098 135300 53104 135312
rect 4028 135272 53104 135300
rect 4028 135260 4034 135272
rect 53098 135260 53104 135272
rect 53156 135260 53162 135312
rect 284202 135260 284208 135312
rect 284260 135300 284266 135312
rect 354674 135300 354680 135312
rect 284260 135272 354680 135300
rect 284260 135260 284266 135272
rect 354674 135260 354680 135272
rect 354732 135260 354738 135312
rect 280893 135235 280951 135241
rect 280893 135201 280905 135235
rect 280939 135232 280951 135235
rect 280982 135232 280988 135244
rect 280939 135204 280988 135232
rect 280939 135201 280951 135204
rect 280893 135195 280951 135201
rect 280982 135192 280988 135204
rect 281040 135192 281046 135244
rect 308490 133900 308496 133952
rect 308548 133940 308554 133952
rect 580166 133940 580172 133952
rect 308548 133912 580172 133940
rect 308548 133900 308554 133912
rect 580166 133900 580172 133912
rect 580224 133900 580230 133952
rect 542354 132472 542360 132524
rect 542412 132512 542418 132524
rect 542630 132512 542636 132524
rect 542412 132484 542636 132512
rect 542412 132472 542418 132484
rect 542630 132472 542636 132484
rect 542688 132472 542694 132524
rect 58526 131112 58532 131164
rect 58584 131152 58590 131164
rect 59354 131152 59360 131164
rect 58584 131124 59360 131152
rect 58584 131112 58590 131124
rect 59354 131112 59360 131124
rect 59412 131112 59418 131164
rect 57238 129752 57244 129804
rect 57296 129792 57302 129804
rect 59722 129792 59728 129804
rect 57296 129764 59728 129792
rect 57296 129752 57302 129764
rect 59722 129752 59728 129764
rect 59780 129752 59786 129804
rect 54754 128324 54760 128376
rect 54812 128364 54818 128376
rect 59354 128364 59360 128376
rect 54812 128336 59360 128364
rect 54812 128324 54818 128336
rect 59354 128324 59360 128336
rect 59412 128324 59418 128376
rect 60642 128324 60648 128376
rect 60700 128364 60706 128376
rect 62390 128364 62396 128376
rect 60700 128336 62396 128364
rect 60700 128324 60706 128336
rect 62390 128324 62396 128336
rect 62448 128324 62454 128376
rect 429286 128324 429292 128376
rect 429344 128364 429350 128376
rect 429470 128364 429476 128376
rect 429344 128336 429476 128364
rect 429344 128324 429350 128336
rect 429470 128324 429476 128336
rect 429528 128324 429534 128376
rect 542354 128256 542360 128308
rect 542412 128296 542418 128308
rect 542630 128296 542636 128308
rect 542412 128268 542636 128296
rect 542412 128256 542418 128268
rect 542630 128256 542636 128268
rect 542688 128256 542694 128308
rect 282178 127576 282184 127628
rect 282236 127616 282242 127628
rect 283558 127616 283564 127628
rect 282236 127588 283564 127616
rect 282236 127576 282242 127588
rect 283558 127576 283564 127588
rect 283616 127576 283622 127628
rect 280890 125712 280896 125724
rect 280851 125684 280896 125712
rect 280890 125672 280896 125684
rect 280948 125672 280954 125724
rect 7929 125579 7987 125585
rect 7929 125545 7941 125579
rect 7975 125576 7987 125579
rect 8018 125576 8024 125588
rect 7975 125548 8024 125576
rect 7975 125545 7987 125548
rect 7929 125539 7987 125545
rect 8018 125536 8024 125548
rect 8076 125536 8082 125588
rect 280890 125576 280896 125588
rect 280851 125548 280896 125576
rect 280890 125536 280896 125548
rect 280948 125536 280954 125588
rect 429286 125576 429292 125588
rect 429247 125548 429292 125576
rect 429286 125536 429292 125548
rect 429344 125536 429350 125588
rect 280798 125468 280804 125520
rect 280856 125508 280862 125520
rect 281350 125508 281356 125520
rect 280856 125480 281356 125508
rect 280856 125468 280862 125480
rect 281350 125468 281356 125480
rect 281408 125468 281414 125520
rect 322290 124108 322296 124160
rect 322348 124148 322354 124160
rect 579890 124148 579896 124160
rect 322348 124120 579896 124148
rect 322348 124108 322354 124120
rect 579890 124108 579896 124120
rect 579948 124108 579954 124160
rect 58434 122884 58440 122936
rect 58492 122924 58498 122936
rect 60274 122924 60280 122936
rect 58492 122896 60280 122924
rect 58492 122884 58498 122896
rect 60274 122884 60280 122896
rect 60332 122884 60338 122936
rect 2774 122136 2780 122188
rect 2832 122176 2838 122188
rect 6178 122176 6184 122188
rect 2832 122148 6184 122176
rect 2832 122136 2838 122148
rect 6178 122136 6184 122148
rect 6236 122136 6242 122188
rect 54662 120096 54668 120148
rect 54720 120136 54726 120148
rect 59354 120136 59360 120148
rect 54720 120108 59360 120136
rect 54720 120096 54726 120108
rect 59354 120096 59360 120108
rect 59412 120096 59418 120148
rect 280798 120096 280804 120148
rect 280856 120136 280862 120148
rect 281166 120136 281172 120148
rect 280856 120108 281172 120136
rect 280856 120096 280862 120108
rect 281166 120096 281172 120108
rect 281224 120096 281230 120148
rect 283834 120096 283840 120148
rect 283892 120136 283898 120148
rect 491294 120136 491300 120148
rect 283892 120108 491300 120136
rect 283892 120096 283898 120108
rect 491294 120096 491300 120108
rect 491352 120096 491358 120148
rect 280890 118640 280896 118652
rect 280851 118612 280896 118640
rect 280890 118600 280896 118612
rect 280948 118600 280954 118652
rect 56042 117308 56048 117360
rect 56100 117348 56106 117360
rect 59354 117348 59360 117360
rect 56100 117320 59360 117348
rect 56100 117308 56106 117320
rect 59354 117308 59360 117320
rect 59412 117308 59418 117360
rect 283650 117308 283656 117360
rect 283708 117348 283714 117360
rect 347866 117348 347872 117360
rect 283708 117320 347872 117348
rect 283708 117308 283714 117320
rect 347866 117308 347872 117320
rect 347924 117308 347930 117360
rect 7926 115988 7932 116000
rect 7887 115960 7932 115988
rect 7926 115948 7932 115960
rect 7984 115948 7990 116000
rect 429286 115988 429292 116000
rect 429247 115960 429292 115988
rect 429286 115948 429292 115960
rect 429344 115948 429350 116000
rect 280893 115923 280951 115929
rect 280893 115889 280905 115923
rect 280939 115920 280951 115923
rect 280982 115920 280988 115932
rect 280939 115892 280988 115920
rect 280939 115889 280951 115892
rect 280893 115883 280951 115889
rect 280982 115880 280988 115892
rect 281040 115880 281046 115932
rect 542354 115880 542360 115932
rect 542412 115920 542418 115932
rect 542538 115920 542544 115932
rect 542412 115892 542544 115920
rect 542412 115880 542418 115892
rect 542538 115880 542544 115892
rect 542596 115880 542602 115932
rect 280798 113908 280804 113960
rect 280856 113948 280862 113960
rect 281166 113948 281172 113960
rect 280856 113920 281172 113948
rect 280856 113908 280862 113920
rect 281166 113908 281172 113920
rect 281224 113908 281230 113960
rect 280798 112344 280804 112396
rect 280856 112384 280862 112396
rect 281350 112384 281356 112396
rect 280856 112356 281356 112384
rect 280856 112344 280862 112356
rect 281350 112344 281356 112356
rect 281408 112344 281414 112396
rect 57146 111800 57152 111852
rect 57204 111840 57210 111852
rect 59630 111840 59636 111852
rect 57204 111812 59636 111840
rect 57204 111800 57210 111812
rect 59630 111800 59636 111812
rect 59688 111800 59694 111852
rect 283742 111800 283748 111852
rect 283800 111840 283806 111852
rect 433334 111840 433340 111852
rect 283800 111812 433340 111840
rect 283800 111800 283806 111812
rect 433334 111800 433340 111812
rect 433392 111800 433398 111852
rect 284018 109012 284024 109064
rect 284076 109052 284082 109064
rect 423674 109052 423680 109064
rect 284076 109024 423680 109052
rect 284076 109012 284082 109024
rect 423674 109012 423680 109024
rect 423732 109012 423738 109064
rect 4062 107652 4068 107704
rect 4120 107692 4126 107704
rect 55766 107692 55772 107704
rect 4120 107664 55772 107692
rect 4120 107652 4126 107664
rect 55766 107652 55772 107664
rect 55824 107652 55830 107704
rect 284018 107652 284024 107704
rect 284076 107692 284082 107704
rect 411254 107692 411260 107704
rect 284076 107664 411260 107692
rect 284076 107652 284082 107664
rect 411254 107652 411260 107664
rect 411312 107652 411318 107704
rect 280798 106496 280804 106548
rect 280856 106536 280862 106548
rect 281350 106536 281356 106548
rect 280856 106508 281356 106536
rect 280856 106496 280862 106508
rect 281350 106496 281356 106508
rect 281408 106496 281414 106548
rect 280890 106332 280896 106344
rect 280851 106304 280896 106332
rect 280890 106292 280896 106304
rect 280948 106292 280954 106344
rect 284018 106292 284024 106344
rect 284076 106332 284082 106344
rect 374086 106332 374092 106344
rect 284076 106304 374092 106332
rect 284076 106292 284082 106304
rect 374086 106292 374092 106304
rect 374144 106292 374150 106344
rect 8018 106264 8024 106276
rect 7979 106236 8024 106264
rect 8018 106224 8024 106236
rect 8076 106224 8082 106276
rect 280798 106224 280804 106276
rect 280856 106264 280862 106276
rect 281166 106264 281172 106276
rect 280856 106236 281172 106264
rect 280856 106224 280862 106236
rect 281166 106224 281172 106236
rect 281224 106224 281230 106276
rect 280890 106196 280896 106208
rect 280851 106168 280896 106196
rect 280890 106156 280896 106168
rect 280948 106156 280954 106208
rect 6178 103504 6184 103556
rect 6236 103544 6242 103556
rect 59354 103544 59360 103556
rect 6236 103516 59360 103544
rect 6236 103504 6242 103516
rect 59354 103504 59360 103516
rect 59412 103504 59418 103556
rect 283834 103504 283840 103556
rect 283892 103544 283898 103556
rect 313274 103544 313280 103556
rect 283892 103516 313280 103544
rect 283892 103504 283898 103516
rect 313274 103504 313280 103516
rect 313332 103504 313338 103556
rect 299658 101436 299664 101448
rect 299619 101408 299664 101436
rect 299658 101396 299664 101408
rect 299716 101396 299722 101448
rect 542630 101436 542636 101448
rect 542591 101408 542636 101436
rect 542630 101396 542636 101408
rect 542688 101396 542694 101448
rect 55950 100716 55956 100768
rect 56008 100756 56014 100768
rect 59354 100756 59360 100768
rect 56008 100728 59360 100756
rect 56008 100716 56014 100728
rect 59354 100716 59360 100728
rect 59412 100716 59418 100768
rect 284202 100716 284208 100768
rect 284260 100756 284266 100768
rect 286226 100756 286232 100768
rect 284260 100728 286232 100756
rect 284260 100716 284266 100728
rect 286226 100716 286232 100728
rect 286284 100716 286290 100768
rect 283650 99356 283656 99408
rect 283708 99396 283714 99408
rect 554038 99396 554044 99408
rect 283708 99368 554044 99396
rect 283708 99356 283714 99368
rect 554038 99356 554044 99368
rect 554096 99356 554102 99408
rect 8018 99328 8024 99340
rect 7979 99300 8024 99328
rect 8018 99288 8024 99300
rect 8076 99288 8082 99340
rect 299658 99328 299664 99340
rect 299619 99300 299664 99328
rect 299658 99288 299664 99300
rect 299716 99288 299722 99340
rect 542633 99331 542691 99337
rect 542633 99297 542645 99331
rect 542679 99328 542691 99331
rect 542722 99328 542728 99340
rect 542679 99300 542728 99328
rect 542679 99297 542691 99300
rect 542633 99291 542691 99297
rect 542722 99288 542728 99300
rect 542780 99288 542786 99340
rect 60090 98880 60096 98932
rect 60148 98920 60154 98932
rect 62298 98920 62304 98932
rect 60148 98892 62304 98920
rect 60148 98880 60154 98892
rect 62298 98880 62304 98892
rect 62356 98880 62362 98932
rect 283834 97996 283840 98048
rect 283892 98036 283898 98048
rect 409138 98036 409144 98048
rect 283892 98008 409144 98036
rect 283892 97996 283898 98008
rect 409138 97996 409144 98008
rect 409196 97996 409202 98048
rect 281074 96840 281080 96892
rect 281132 96840 281138 96892
rect 281092 96688 281120 96840
rect 280893 96679 280951 96685
rect 280893 96645 280905 96679
rect 280939 96676 280951 96679
rect 280982 96676 280988 96688
rect 280939 96648 280988 96676
rect 280939 96645 280951 96648
rect 280893 96639 280951 96645
rect 280982 96636 280988 96648
rect 281040 96636 281046 96688
rect 281074 96636 281080 96688
rect 281132 96636 281138 96688
rect 429102 96568 429108 96620
rect 429160 96608 429166 96620
rect 429378 96608 429384 96620
rect 429160 96580 429384 96608
rect 429160 96568 429166 96580
rect 429378 96568 429384 96580
rect 429436 96568 429442 96620
rect 280982 96540 280988 96552
rect 280943 96512 280988 96540
rect 280982 96500 280988 96512
rect 281040 96500 281046 96552
rect 283834 95208 283840 95260
rect 283892 95248 283898 95260
rect 389818 95248 389824 95260
rect 283892 95220 389824 95248
rect 283892 95208 283898 95220
rect 389818 95208 389824 95220
rect 389876 95208 389882 95260
rect 280798 94596 280804 94648
rect 280856 94636 280862 94648
rect 281166 94636 281172 94648
rect 280856 94608 281172 94636
rect 280856 94596 280862 94608
rect 281166 94596 281172 94608
rect 281224 94596 281230 94648
rect 280798 94460 280804 94512
rect 280856 94500 280862 94512
rect 281350 94500 281356 94512
rect 280856 94472 281356 94500
rect 280856 94460 280862 94472
rect 281350 94460 281356 94472
rect 281408 94460 281414 94512
rect 283834 93780 283840 93832
rect 283892 93820 283898 93832
rect 290458 93820 290464 93832
rect 283892 93792 290464 93820
rect 283892 93780 283898 93792
rect 290458 93780 290464 93792
rect 290516 93780 290522 93832
rect 8110 90992 8116 91044
rect 8168 91032 8174 91044
rect 59354 91032 59360 91044
rect 8168 91004 59360 91032
rect 8168 90992 8174 91004
rect 59354 90992 59360 91004
rect 59412 90992 59418 91044
rect 284018 89700 284024 89752
rect 284076 89740 284082 89752
rect 469214 89740 469220 89752
rect 284076 89712 469220 89740
rect 284076 89700 284082 89712
rect 469214 89700 469220 89712
rect 469272 89700 469278 89752
rect 280982 89672 280988 89684
rect 280943 89644 280988 89672
rect 280982 89632 280988 89644
rect 281040 89632 281046 89684
rect 283834 89632 283840 89684
rect 283892 89672 283898 89684
rect 308490 89672 308496 89684
rect 283892 89644 308496 89672
rect 283892 89632 283898 89644
rect 308490 89632 308496 89644
rect 308548 89632 308554 89684
rect 501598 88272 501604 88324
rect 501656 88312 501662 88324
rect 579890 88312 579896 88324
rect 501656 88284 579896 88312
rect 501656 88272 501662 88284
rect 579890 88272 579896 88284
rect 579948 88272 579954 88324
rect 283834 86980 283840 87032
rect 283892 87020 283898 87032
rect 318058 87020 318064 87032
rect 283892 86992 318064 87020
rect 283892 86980 283898 86992
rect 318058 86980 318064 86992
rect 318116 86980 318122 87032
rect 280893 86955 280951 86961
rect 280893 86921 280905 86955
rect 280939 86952 280951 86955
rect 280982 86952 280988 86964
rect 280939 86924 280988 86952
rect 280939 86921 280951 86924
rect 280893 86915 280951 86921
rect 280982 86912 280988 86924
rect 281040 86912 281046 86964
rect 299658 86952 299664 86964
rect 299619 86924 299664 86952
rect 299658 86912 299664 86924
rect 299716 86912 299722 86964
rect 287882 86232 287888 86284
rect 287940 86272 287946 86284
rect 331306 86272 331312 86284
rect 287940 86244 331312 86272
rect 287940 86232 287946 86244
rect 331306 86232 331312 86244
rect 331364 86232 331370 86284
rect 283834 85552 283840 85604
rect 283892 85592 283898 85604
rect 433426 85592 433432 85604
rect 283892 85564 433432 85592
rect 283892 85552 283898 85564
rect 433426 85552 433432 85564
rect 433484 85552 433490 85604
rect 280798 85008 280804 85060
rect 280856 85048 280862 85060
rect 281442 85048 281448 85060
rect 280856 85020 281448 85048
rect 280856 85008 280862 85020
rect 281442 85008 281448 85020
rect 281500 85008 281506 85060
rect 280798 84872 280804 84924
rect 280856 84912 280862 84924
rect 281350 84912 281356 84924
rect 280856 84884 281356 84912
rect 280856 84872 280862 84884
rect 281350 84872 281356 84884
rect 281408 84872 281414 84924
rect 283650 81404 283656 81456
rect 283708 81444 283714 81456
rect 286502 81444 286508 81456
rect 283708 81416 286508 81444
rect 283708 81404 283714 81416
rect 286502 81404 286508 81416
rect 286560 81404 286566 81456
rect 429286 80044 429292 80096
rect 429344 80044 429350 80096
rect 3970 79976 3976 80028
rect 4028 80016 4034 80028
rect 55858 80016 55864 80028
rect 4028 79988 55864 80016
rect 4028 79976 4034 79988
rect 55858 79976 55864 79988
rect 55916 79976 55922 80028
rect 429304 79948 429332 80044
rect 429378 79948 429384 79960
rect 429304 79920 429384 79948
rect 429378 79908 429384 79920
rect 429436 79908 429442 79960
rect 284202 78684 284208 78736
rect 284260 78724 284266 78736
rect 403618 78724 403624 78736
rect 284260 78696 403624 78724
rect 284260 78684 284266 78696
rect 403618 78684 403624 78696
rect 403676 78684 403682 78736
rect 10318 78616 10324 78668
rect 10376 78656 10382 78668
rect 59354 78656 59360 78668
rect 10376 78628 59360 78656
rect 10376 78616 10382 78628
rect 59354 78616 59360 78628
rect 59412 78616 59418 78668
rect 280890 77296 280896 77308
rect 280851 77268 280896 77296
rect 280890 77256 280896 77268
rect 280948 77256 280954 77308
rect 299658 77296 299664 77308
rect 299619 77268 299664 77296
rect 299658 77256 299664 77268
rect 299716 77256 299722 77308
rect 62206 77228 62212 77240
rect 62167 77200 62212 77228
rect 62206 77188 62212 77200
rect 62264 77188 62270 77240
rect 280982 77228 280988 77240
rect 280943 77200 280988 77228
rect 280982 77188 280988 77200
rect 281040 77188 281046 77240
rect 294690 77188 294696 77240
rect 294748 77228 294754 77240
rect 579614 77228 579620 77240
rect 294748 77200 579620 77228
rect 294748 77188 294754 77200
rect 579614 77188 579620 77200
rect 579672 77188 579678 77240
rect 280798 75284 280804 75336
rect 280856 75324 280862 75336
rect 281350 75324 281356 75336
rect 280856 75296 281356 75324
rect 280856 75284 280862 75296
rect 281350 75284 281356 75296
rect 281408 75284 281414 75336
rect 280798 75148 280804 75200
rect 280856 75188 280862 75200
rect 281442 75188 281448 75200
rect 280856 75160 281448 75188
rect 280856 75148 280862 75160
rect 281442 75148 281448 75160
rect 281500 75148 281506 75200
rect 55858 74536 55864 74588
rect 55916 74576 55922 74588
rect 59354 74576 59360 74588
rect 55916 74548 59360 74576
rect 55916 74536 55922 74548
rect 59354 74536 59360 74548
rect 59412 74536 59418 74588
rect 284202 74536 284208 74588
rect 284260 74576 284266 74588
rect 358814 74576 358820 74588
rect 284260 74548 358820 74576
rect 284260 74536 284266 74548
rect 358814 74536 358820 74548
rect 358872 74536 358878 74588
rect 284202 71748 284208 71800
rect 284260 71788 284266 71800
rect 334618 71788 334624 71800
rect 284260 71760 334624 71788
rect 284260 71748 284266 71760
rect 334618 71748 334624 71760
rect 334676 71748 334682 71800
rect 280890 67668 280896 67720
rect 280948 67708 280954 67720
rect 280985 67711 281043 67717
rect 280985 67708 280997 67711
rect 280948 67680 280997 67708
rect 280948 67668 280954 67680
rect 280985 67677 280997 67680
rect 281031 67677 281043 67711
rect 280985 67671 281043 67677
rect 62209 67643 62267 67649
rect 62209 67609 62221 67643
rect 62255 67640 62267 67643
rect 62298 67640 62304 67652
rect 62255 67612 62304 67640
rect 62255 67609 62267 67612
rect 62209 67603 62267 67609
rect 62298 67600 62304 67612
rect 62356 67600 62362 67652
rect 283834 67600 283840 67652
rect 283892 67640 283898 67652
rect 496078 67640 496084 67652
rect 283892 67612 496084 67640
rect 283892 67600 283898 67612
rect 496078 67600 496084 67612
rect 496136 67600 496142 67652
rect 280890 67572 280896 67584
rect 280851 67544 280896 67572
rect 280890 67532 280896 67544
rect 280948 67532 280954 67584
rect 299658 67572 299664 67584
rect 299619 67544 299664 67572
rect 299658 67532 299664 67544
rect 299716 67532 299722 67584
rect 542538 67532 542544 67584
rect 542596 67572 542602 67584
rect 542722 67572 542728 67584
rect 542596 67544 542728 67572
rect 542596 67532 542602 67544
rect 542722 67532 542728 67544
rect 542780 67532 542786 67584
rect 280798 67396 280804 67448
rect 280856 67436 280862 67448
rect 281442 67436 281448 67448
rect 280856 67408 281448 67436
rect 280856 67396 280862 67408
rect 281442 67396 281448 67408
rect 281500 67396 281506 67448
rect 280798 65424 280804 65476
rect 280856 65464 280862 65476
rect 281350 65464 281356 65476
rect 280856 65436 281356 65464
rect 280856 65424 280862 65436
rect 281350 65424 281356 65436
rect 281408 65424 281414 65476
rect 55674 65288 55680 65340
rect 55732 65328 55738 65340
rect 59354 65328 59360 65340
rect 55732 65300 59360 65328
rect 55732 65288 55738 65300
rect 59354 65288 59360 65300
rect 59412 65288 59418 65340
rect 407758 64812 407764 64864
rect 407816 64852 407822 64864
rect 580166 64852 580172 64864
rect 407816 64824 580172 64852
rect 407816 64812 407822 64824
rect 580166 64812 580172 64824
rect 580224 64812 580230 64864
rect 283834 63520 283840 63572
rect 283892 63560 283898 63572
rect 289906 63560 289912 63572
rect 283892 63532 289912 63560
rect 283892 63520 283898 63532
rect 289906 63520 289912 63532
rect 289964 63520 289970 63572
rect 283834 62024 283840 62076
rect 283892 62064 283898 62076
rect 304350 62064 304356 62076
rect 283892 62036 304356 62064
rect 283892 62024 283898 62036
rect 304350 62024 304356 62036
rect 304408 62024 304414 62076
rect 299658 60976 299664 60988
rect 299619 60948 299664 60976
rect 299658 60936 299664 60948
rect 299716 60936 299722 60988
rect 4798 60664 4804 60716
rect 4856 60704 4862 60716
rect 59354 60704 59360 60716
rect 4856 60676 59360 60704
rect 4856 60664 4862 60676
rect 59354 60664 59360 60676
rect 59412 60664 59418 60716
rect 280893 60639 280951 60645
rect 280893 60605 280905 60639
rect 280939 60636 280951 60639
rect 280982 60636 280988 60648
rect 280939 60608 280988 60636
rect 280939 60605 280951 60608
rect 280893 60599 280951 60605
rect 280982 60596 280988 60608
rect 281040 60596 281046 60648
rect 429378 60596 429384 60648
rect 429436 60636 429442 60648
rect 429562 60636 429568 60648
rect 429436 60608 429568 60636
rect 429436 60596 429442 60608
rect 429562 60596 429568 60608
rect 429620 60596 429626 60648
rect 283834 57944 283840 57996
rect 283892 57984 283898 57996
rect 494698 57984 494704 57996
rect 283892 57956 494704 57984
rect 283892 57944 283898 57956
rect 494698 57944 494704 57956
rect 494756 57944 494762 57996
rect 280893 52751 280951 52757
rect 280893 52717 280905 52751
rect 280939 52748 280951 52751
rect 281350 52748 281356 52760
rect 280939 52720 281356 52748
rect 280939 52717 280951 52720
rect 280893 52711 280951 52717
rect 281350 52708 281356 52720
rect 281408 52708 281414 52760
rect 337378 51688 337384 51740
rect 337436 51728 337442 51740
rect 538214 51728 538220 51740
rect 337436 51700 538220 51728
rect 337436 51688 337442 51700
rect 538214 51688 538220 51700
rect 538272 51688 538278 51740
rect 281442 51116 281448 51128
rect 280816 51088 281448 51116
rect 280816 51060 280844 51088
rect 281442 51076 281448 51088
rect 281500 51076 281506 51128
rect 280798 51008 280804 51060
rect 280856 51008 280862 51060
rect 280982 51008 280988 51060
rect 281040 51048 281046 51060
rect 281350 51048 281356 51060
rect 281040 51020 281356 51048
rect 281040 51008 281046 51020
rect 281350 51008 281356 51020
rect 281408 51008 281414 51060
rect 305638 50328 305644 50380
rect 305696 50368 305702 50380
rect 459646 50368 459652 50380
rect 305696 50340 459652 50368
rect 305696 50328 305702 50340
rect 459646 50328 459652 50340
rect 459704 50328 459710 50380
rect 280890 48328 280896 48340
rect 280851 48300 280896 48328
rect 280890 48288 280896 48300
rect 280948 48288 280954 48340
rect 280798 48220 280804 48272
rect 280856 48260 280862 48272
rect 281350 48260 281356 48272
rect 280856 48232 281356 48260
rect 280856 48220 280862 48232
rect 281350 48220 281356 48232
rect 281408 48220 281414 48272
rect 318058 47540 318064 47592
rect 318116 47580 318122 47592
rect 561674 47580 561680 47592
rect 318116 47552 561680 47580
rect 318116 47540 318122 47552
rect 561674 47540 561680 47552
rect 561732 47540 561738 47592
rect 283834 45568 283840 45620
rect 283892 45608 283898 45620
rect 386414 45608 386420 45620
rect 283892 45580 386420 45608
rect 283892 45568 283898 45580
rect 386414 45568 386420 45580
rect 386472 45568 386478 45620
rect 287790 44820 287796 44872
rect 287848 44860 287854 44872
rect 310514 44860 310520 44872
rect 287848 44832 310520 44860
rect 287848 44820 287854 44832
rect 310514 44820 310520 44832
rect 310572 44820 310578 44872
rect 62206 44276 62212 44328
rect 62264 44316 62270 44328
rect 62264 44288 277072 44316
rect 62264 44276 62270 44288
rect 277044 43920 277072 44288
rect 283834 44140 283840 44192
rect 283892 44180 283898 44192
rect 506474 44180 506480 44192
rect 283892 44152 506480 44180
rect 283892 44140 283898 44152
rect 506474 44140 506480 44152
rect 506532 44140 506538 44192
rect 277026 43868 277032 43920
rect 277084 43868 277090 43920
rect 60458 43800 60464 43852
rect 60516 43840 60522 43852
rect 144178 43840 144184 43852
rect 60516 43812 144184 43840
rect 60516 43800 60522 43812
rect 144178 43800 144184 43812
rect 144236 43800 144242 43852
rect 61010 43732 61016 43784
rect 61068 43772 61074 43784
rect 149057 43775 149115 43781
rect 149057 43772 149069 43775
rect 61068 43744 149069 43772
rect 61068 43732 61074 43744
rect 149057 43741 149069 43744
rect 149103 43741 149115 43775
rect 149057 43735 149115 43741
rect 61286 43664 61292 43716
rect 61344 43704 61350 43716
rect 187694 43704 187700 43716
rect 61344 43676 187700 43704
rect 61344 43664 61350 43676
rect 187694 43664 187700 43676
rect 187752 43664 187758 43716
rect 211062 43664 211068 43716
rect 211120 43704 211126 43716
rect 283098 43704 283104 43716
rect 211120 43676 283104 43704
rect 211120 43664 211126 43676
rect 283098 43664 283104 43676
rect 283156 43664 283162 43716
rect 62022 43596 62028 43648
rect 62080 43636 62086 43648
rect 223850 43636 223856 43648
rect 62080 43608 223856 43636
rect 62080 43596 62086 43608
rect 223850 43596 223856 43608
rect 223908 43596 223914 43648
rect 59998 43528 60004 43580
rect 60056 43568 60062 43580
rect 227714 43568 227720 43580
rect 60056 43540 227720 43568
rect 60056 43528 60062 43540
rect 227714 43528 227720 43540
rect 227772 43528 227778 43580
rect 60274 43460 60280 43512
rect 60332 43500 60338 43512
rect 333974 43500 333980 43512
rect 60332 43472 333980 43500
rect 60332 43460 60338 43472
rect 333974 43460 333980 43472
rect 334032 43460 334038 43512
rect 334618 43460 334624 43512
rect 334676 43500 334682 43512
rect 534074 43500 534080 43512
rect 334676 43472 534080 43500
rect 334676 43460 334682 43472
rect 534074 43460 534080 43472
rect 534132 43460 534138 43512
rect 3418 43392 3424 43444
rect 3476 43432 3482 43444
rect 57054 43432 57060 43444
rect 3476 43404 57060 43432
rect 3476 43392 3482 43404
rect 57054 43392 57060 43404
rect 57112 43392 57118 43444
rect 61470 43392 61476 43444
rect 61528 43432 61534 43444
rect 362954 43432 362960 43444
rect 61528 43404 362960 43432
rect 61528 43392 61534 43404
rect 362954 43392 362960 43404
rect 363012 43392 363018 43444
rect 60366 42916 60372 42968
rect 60424 42956 60430 42968
rect 64138 42956 64144 42968
rect 60424 42928 64144 42956
rect 60424 42916 60430 42928
rect 64138 42916 64144 42928
rect 64196 42916 64202 42968
rect 200022 42848 200028 42900
rect 200080 42888 200086 42900
rect 286318 42888 286324 42900
rect 200080 42860 286324 42888
rect 200080 42848 200086 42860
rect 286318 42848 286324 42860
rect 286376 42848 286382 42900
rect 233510 42780 233516 42832
rect 233568 42820 233574 42832
rect 429378 42820 429384 42832
rect 233568 42792 429384 42820
rect 233568 42780 233574 42792
rect 429378 42780 429384 42792
rect 429436 42780 429442 42832
rect 248414 42712 248420 42764
rect 248472 42752 248478 42764
rect 286410 42752 286416 42764
rect 248472 42724 286416 42752
rect 248472 42712 248478 42724
rect 286410 42712 286416 42724
rect 286468 42712 286474 42764
rect 94222 42644 94228 42696
rect 94280 42684 94286 42696
rect 285122 42684 285128 42696
rect 94280 42656 285128 42684
rect 94280 42644 94286 42656
rect 285122 42644 285128 42656
rect 285180 42644 285186 42696
rect 55766 42576 55772 42628
rect 55824 42616 55830 42628
rect 160462 42616 160468 42628
rect 55824 42588 160468 42616
rect 55824 42576 55830 42588
rect 160462 42576 160468 42588
rect 160520 42576 160526 42628
rect 185118 42576 185124 42628
rect 185176 42616 185182 42628
rect 290550 42616 290556 42628
rect 185176 42588 290556 42616
rect 185176 42576 185182 42588
rect 290550 42576 290556 42588
rect 290608 42576 290614 42628
rect 53098 42508 53104 42560
rect 53156 42548 53162 42560
rect 146478 42548 146484 42560
rect 53156 42520 146484 42548
rect 53156 42508 53162 42520
rect 146478 42508 146484 42520
rect 146536 42508 146542 42560
rect 191006 42508 191012 42560
rect 191064 42548 191070 42560
rect 291930 42548 291936 42560
rect 191064 42520 291936 42548
rect 191064 42508 191070 42520
rect 291930 42508 291936 42520
rect 291988 42508 291994 42560
rect 195054 42440 195060 42492
rect 195112 42480 195118 42492
rect 287698 42480 287704 42492
rect 195112 42452 287704 42480
rect 195112 42440 195118 42452
rect 287698 42440 287704 42452
rect 287756 42440 287762 42492
rect 168282 42372 168288 42424
rect 168340 42412 168346 42424
rect 286134 42412 286140 42424
rect 168340 42384 286140 42412
rect 168340 42372 168346 42384
rect 286134 42372 286140 42384
rect 286192 42372 286198 42424
rect 157242 42304 157248 42356
rect 157300 42344 157306 42356
rect 286226 42344 286232 42356
rect 157300 42316 286232 42344
rect 157300 42304 157306 42316
rect 286226 42304 286232 42316
rect 286284 42304 286290 42356
rect 41322 42236 41328 42288
rect 41380 42276 41386 42288
rect 96522 42276 96528 42288
rect 41380 42248 96528 42276
rect 41380 42236 41386 42248
rect 96522 42236 96528 42248
rect 96580 42236 96586 42288
rect 155862 42236 155868 42288
rect 155920 42276 155926 42288
rect 287238 42276 287244 42288
rect 155920 42248 287244 42276
rect 155920 42236 155926 42248
rect 287238 42236 287244 42248
rect 287296 42236 287302 42288
rect 56226 42168 56232 42220
rect 56284 42208 56290 42220
rect 137005 42211 137063 42217
rect 137005 42208 137017 42211
rect 56284 42180 137017 42208
rect 56284 42168 56290 42180
rect 137005 42177 137017 42180
rect 137051 42177 137063 42211
rect 137005 42171 137063 42177
rect 154482 42168 154488 42220
rect 154540 42208 154546 42220
rect 285950 42208 285956 42220
rect 154540 42180 285956 42208
rect 154540 42168 154546 42180
rect 285950 42168 285956 42180
rect 286008 42168 286014 42220
rect 56318 42100 56324 42152
rect 56376 42140 56382 42152
rect 128446 42140 128452 42152
rect 56376 42112 128452 42140
rect 56376 42100 56382 42112
rect 128446 42100 128452 42112
rect 128504 42100 128510 42152
rect 135073 42143 135131 42149
rect 135073 42109 135085 42143
rect 135119 42140 135131 42143
rect 286042 42140 286048 42152
rect 135119 42112 286048 42140
rect 135119 42109 135131 42112
rect 135073 42103 135131 42109
rect 286042 42100 286048 42112
rect 286100 42100 286106 42152
rect 3510 42032 3516 42084
rect 3568 42072 3574 42084
rect 88978 42072 88984 42084
rect 3568 42044 88984 42072
rect 3568 42032 3574 42044
rect 88978 42032 88984 42044
rect 89036 42032 89042 42084
rect 128354 42032 128360 42084
rect 128412 42072 128418 42084
rect 580258 42072 580264 42084
rect 128412 42044 580264 42072
rect 128412 42032 128418 42044
rect 580258 42032 580264 42044
rect 580316 42032 580322 42084
rect 255406 41964 255412 42016
rect 255464 42004 255470 42016
rect 285306 42004 285312 42016
rect 255464 41976 285312 42004
rect 255464 41964 255470 41976
rect 285306 41964 285312 41976
rect 285364 41964 285370 42016
rect 51718 41896 51724 41948
rect 51776 41936 51782 41948
rect 258350 41936 258356 41948
rect 51776 41908 258356 41936
rect 51776 41896 51782 41908
rect 258350 41896 258356 41908
rect 258408 41896 258414 41948
rect 262122 41896 262128 41948
rect 262180 41936 262186 41948
rect 288710 41936 288716 41948
rect 262180 41908 288716 41936
rect 262180 41896 262186 41908
rect 288710 41896 288716 41908
rect 288768 41896 288774 41948
rect 279418 41420 279424 41472
rect 279476 41460 279482 41472
rect 284662 41460 284668 41472
rect 279476 41432 284668 41460
rect 279476 41420 279482 41432
rect 284662 41420 284668 41432
rect 284720 41420 284726 41472
rect 8938 41352 8944 41404
rect 8996 41392 9002 41404
rect 88150 41392 88156 41404
rect 8996 41364 88156 41392
rect 8996 41352 9002 41364
rect 88150 41352 88156 41364
rect 88208 41352 88214 41404
rect 96522 41352 96528 41404
rect 96580 41392 96586 41404
rect 216766 41392 216772 41404
rect 96580 41364 216772 41392
rect 96580 41352 96586 41364
rect 216766 41352 216772 41364
rect 216824 41352 216830 41404
rect 494698 41352 494704 41404
rect 494756 41392 494762 41404
rect 580166 41392 580172 41404
rect 494756 41364 580172 41392
rect 494756 41352 494762 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 7558 41284 7564 41336
rect 7616 41324 7622 41336
rect 127710 41324 127716 41336
rect 7616 41296 127716 41324
rect 7616 41284 7622 41296
rect 127710 41284 127716 41296
rect 127768 41284 127774 41336
rect 137002 41324 137008 41336
rect 136963 41296 137008 41324
rect 137002 41284 137008 41296
rect 137060 41284 137066 41336
rect 270126 41284 270132 41336
rect 270184 41324 270190 41336
rect 338114 41324 338120 41336
rect 270184 41296 338120 41324
rect 270184 41284 270190 41296
rect 338114 41284 338120 41296
rect 338172 41284 338178 41336
rect 88978 41216 88984 41268
rect 89036 41256 89042 41268
rect 97166 41256 97172 41268
rect 89036 41228 97172 41256
rect 89036 41216 89042 41228
rect 97166 41216 97172 41228
rect 97224 41216 97230 41268
rect 105998 41216 106004 41268
rect 106056 41256 106062 41268
rect 128354 41256 128360 41268
rect 106056 41228 128360 41256
rect 106056 41216 106062 41228
rect 128354 41216 128360 41228
rect 128412 41216 128418 41268
rect 181254 41216 181260 41268
rect 181312 41256 181318 41268
rect 182082 41256 182088 41268
rect 181312 41228 182088 41256
rect 181312 41216 181318 41228
rect 182082 41216 182088 41228
rect 182140 41216 182146 41268
rect 210878 41256 210884 41268
rect 205008 41228 210884 41256
rect 57054 41148 57060 41200
rect 57112 41188 57118 41200
rect 143534 41188 143540 41200
rect 57112 41160 143540 41188
rect 57112 41148 57118 41160
rect 143534 41148 143540 41160
rect 143592 41148 143598 41200
rect 197998 41148 198004 41200
rect 198056 41188 198062 41200
rect 204898 41188 204904 41200
rect 198056 41160 204904 41188
rect 198056 41148 198062 41160
rect 204898 41148 204904 41160
rect 204956 41148 204962 41200
rect 11698 41080 11704 41132
rect 11756 41120 11762 41132
rect 89254 41120 89260 41132
rect 11756 41092 89260 41120
rect 11756 41080 11762 41092
rect 89254 41080 89260 41092
rect 89312 41080 89318 41132
rect 103974 41080 103980 41132
rect 104032 41120 104038 41132
rect 121454 41120 121460 41132
rect 104032 41092 121460 41120
rect 104032 41080 104038 41092
rect 121454 41080 121460 41092
rect 121512 41080 121518 41132
rect 158622 41080 158628 41132
rect 158680 41120 158686 41132
rect 205008 41120 205036 41228
rect 210878 41216 210884 41228
rect 210936 41216 210942 41268
rect 229646 41216 229652 41268
rect 229704 41256 229710 41268
rect 239398 41256 239404 41268
rect 229704 41228 239404 41256
rect 229704 41216 229710 41228
rect 239398 41216 239404 41228
rect 239456 41216 239462 41268
rect 257246 41216 257252 41268
rect 257304 41256 257310 41268
rect 365714 41256 365720 41268
rect 257304 41228 365720 41256
rect 257304 41216 257310 41228
rect 365714 41216 365720 41228
rect 365772 41216 365778 41268
rect 208302 41148 208308 41200
rect 208360 41188 208366 41200
rect 211798 41188 211804 41200
rect 208360 41160 211804 41188
rect 208360 41148 208366 41160
rect 211798 41148 211804 41160
rect 211856 41148 211862 41200
rect 239582 41148 239588 41200
rect 239640 41188 239646 41200
rect 380894 41188 380900 41200
rect 239640 41160 380900 41188
rect 239640 41148 239646 41160
rect 380894 41148 380900 41160
rect 380952 41148 380958 41200
rect 158680 41092 205036 41120
rect 158680 41080 158686 41092
rect 234614 41080 234620 41132
rect 234672 41120 234678 41132
rect 405734 41120 405740 41132
rect 234672 41092 405740 41120
rect 234672 41080 234678 41092
rect 405734 41080 405740 41092
rect 405792 41080 405798 41132
rect 3602 41012 3608 41064
rect 3660 41052 3666 41064
rect 106918 41052 106924 41064
rect 3660 41024 106924 41052
rect 3660 41012 3666 41024
rect 106918 41012 106924 41024
rect 106976 41012 106982 41064
rect 139670 41012 139676 41064
rect 139728 41052 139734 41064
rect 356054 41052 356060 41064
rect 139728 41024 356060 41052
rect 139728 41012 139734 41024
rect 356054 41012 356060 41024
rect 356112 41012 356118 41064
rect 128814 40944 128820 40996
rect 128872 40984 128878 40996
rect 129642 40984 129648 40996
rect 128872 40956 129648 40984
rect 128872 40944 128878 40956
rect 129642 40944 129648 40956
rect 129700 40944 129706 40996
rect 153470 40944 153476 40996
rect 153528 40984 153534 40996
rect 383654 40984 383660 40996
rect 153528 40956 383660 40984
rect 153528 40944 153534 40956
rect 383654 40944 383660 40956
rect 383712 40944 383718 40996
rect 2682 40876 2688 40928
rect 2740 40916 2746 40928
rect 235534 40916 235540 40928
rect 2740 40888 235540 40916
rect 2740 40876 2746 40888
rect 235534 40876 235540 40888
rect 235592 40876 235598 40928
rect 245470 40876 245476 40928
rect 245528 40916 245534 40928
rect 441614 40916 441620 40928
rect 245528 40888 441620 40916
rect 245528 40876 245534 40888
rect 441614 40876 441620 40888
rect 441672 40876 441678 40928
rect 87230 40808 87236 40860
rect 87288 40848 87294 40860
rect 322934 40848 322940 40860
rect 87288 40820 322940 40848
rect 87288 40808 87294 40820
rect 322934 40808 322940 40820
rect 322992 40808 322998 40860
rect 83182 40740 83188 40792
rect 83240 40780 83246 40792
rect 115198 40780 115204 40792
rect 83240 40752 115204 40780
rect 83240 40740 83246 40752
rect 115198 40740 115204 40752
rect 115256 40740 115262 40792
rect 164326 40740 164332 40792
rect 164384 40780 164390 40792
rect 407758 40780 407764 40792
rect 164384 40752 407764 40780
rect 164384 40740 164390 40752
rect 407758 40740 407764 40752
rect 407816 40740 407822 40792
rect 111886 40672 111892 40724
rect 111944 40712 111950 40724
rect 376754 40712 376760 40724
rect 111944 40684 376760 40712
rect 111944 40672 111950 40684
rect 376754 40672 376760 40684
rect 376812 40672 376818 40724
rect 240502 40196 240508 40248
rect 240560 40236 240566 40248
rect 241238 40236 241244 40248
rect 240560 40208 241244 40236
rect 240560 40196 240566 40208
rect 241238 40196 241244 40208
rect 241296 40196 241302 40248
rect 249334 40128 249340 40180
rect 249392 40168 249398 40180
rect 255958 40168 255964 40180
rect 249392 40140 255964 40168
rect 249392 40128 249398 40140
rect 255958 40128 255964 40140
rect 256016 40128 256022 40180
rect 63494 40060 63500 40112
rect 63552 40100 63558 40112
rect 65518 40100 65524 40112
rect 63552 40072 65524 40100
rect 63552 40060 63558 40072
rect 65518 40060 65524 40072
rect 65576 40060 65582 40112
rect 69382 40060 69388 40112
rect 69440 40100 69446 40112
rect 70302 40100 70308 40112
rect 69440 40072 70308 40100
rect 69440 40060 69446 40072
rect 70302 40060 70308 40072
rect 70360 40060 70366 40112
rect 70486 40060 70492 40112
rect 70544 40100 70550 40112
rect 71682 40100 71688 40112
rect 70544 40072 71688 40100
rect 70544 40060 70550 40072
rect 71682 40060 71688 40072
rect 71740 40060 71746 40112
rect 84286 40060 84292 40112
rect 84344 40100 84350 40112
rect 85482 40100 85488 40112
rect 84344 40072 85488 40100
rect 84344 40060 84350 40072
rect 85482 40060 85488 40072
rect 85540 40060 85546 40112
rect 91094 40060 91100 40112
rect 91152 40100 91158 40112
rect 92290 40100 92296 40112
rect 91152 40072 92296 40100
rect 91152 40060 91158 40072
rect 92290 40060 92296 40072
rect 92348 40060 92354 40112
rect 110966 40060 110972 40112
rect 111024 40100 111030 40112
rect 111702 40100 111708 40112
rect 111024 40072 111708 40100
rect 111024 40060 111030 40072
rect 111702 40060 111708 40072
rect 111760 40060 111766 40112
rect 114830 40060 114836 40112
rect 114888 40100 114894 40112
rect 115842 40100 115848 40112
rect 114888 40072 115848 40100
rect 114888 40060 114894 40072
rect 115842 40060 115848 40072
rect 115900 40060 115906 40112
rect 118878 40060 118884 40112
rect 118936 40100 118942 40112
rect 119890 40100 119896 40112
rect 118936 40072 119896 40100
rect 118936 40060 118942 40072
rect 119890 40060 119896 40072
rect 119948 40060 119954 40112
rect 125870 40060 125876 40112
rect 125928 40100 125934 40112
rect 126790 40100 126796 40112
rect 125928 40072 126796 40100
rect 125928 40060 125934 40072
rect 126790 40060 126796 40072
rect 126848 40060 126854 40112
rect 129734 40060 129740 40112
rect 129792 40100 129798 40112
rect 131022 40100 131028 40112
rect 129792 40072 131028 40100
rect 129792 40060 129798 40072
rect 131022 40060 131028 40072
rect 131080 40060 131086 40112
rect 132678 40060 132684 40112
rect 132736 40100 132742 40112
rect 133782 40100 133788 40112
rect 132736 40072 133788 40100
rect 132736 40060 132742 40072
rect 133782 40060 133788 40072
rect 133840 40060 133846 40112
rect 135622 40060 135628 40112
rect 135680 40100 135686 40112
rect 136450 40100 136456 40112
rect 135680 40072 136456 40100
rect 135680 40060 135686 40072
rect 136450 40060 136456 40072
rect 136508 40060 136514 40112
rect 136726 40060 136732 40112
rect 136784 40100 136790 40112
rect 137922 40100 137928 40112
rect 136784 40072 137928 40100
rect 136784 40060 136790 40072
rect 137922 40060 137928 40072
rect 137980 40060 137986 40112
rect 142614 40060 142620 40112
rect 142672 40100 142678 40112
rect 143442 40100 143448 40112
rect 142672 40072 143448 40100
rect 142672 40060 142678 40072
rect 143442 40060 143448 40072
rect 143500 40060 143506 40112
rect 149606 40060 149612 40112
rect 149664 40100 149670 40112
rect 150342 40100 150348 40112
rect 149664 40072 150348 40100
rect 149664 40060 149670 40072
rect 150342 40060 150348 40072
rect 150400 40060 150406 40112
rect 157518 40060 157524 40112
rect 157576 40100 157582 40112
rect 158530 40100 158536 40112
rect 157576 40072 158536 40100
rect 157576 40060 157582 40072
rect 158530 40060 158536 40072
rect 158588 40060 158594 40112
rect 163406 40060 163412 40112
rect 163464 40100 163470 40112
rect 164142 40100 164148 40112
rect 163464 40072 164148 40100
rect 163464 40060 163470 40072
rect 164142 40060 164148 40072
rect 164200 40060 164206 40112
rect 167270 40060 167276 40112
rect 167328 40100 167334 40112
rect 168190 40100 168196 40112
rect 167328 40072 168196 40100
rect 167328 40060 167334 40072
rect 168190 40060 168196 40072
rect 168248 40060 168254 40112
rect 170214 40060 170220 40112
rect 170272 40100 170278 40112
rect 171042 40100 171048 40112
rect 170272 40072 171048 40100
rect 170272 40060 170278 40072
rect 171042 40060 171048 40072
rect 171100 40060 171106 40112
rect 171318 40060 171324 40112
rect 171376 40100 171382 40112
rect 172330 40100 172336 40112
rect 171376 40072 172336 40100
rect 171376 40060 171382 40072
rect 172330 40060 172336 40072
rect 172388 40060 172394 40112
rect 174262 40060 174268 40112
rect 174320 40100 174326 40112
rect 175182 40100 175188 40112
rect 174320 40072 175188 40100
rect 174320 40060 174326 40072
rect 175182 40060 175188 40072
rect 175240 40060 175246 40112
rect 178126 40060 178132 40112
rect 178184 40100 178190 40112
rect 179230 40100 179236 40112
rect 178184 40072 179236 40100
rect 178184 40060 178190 40072
rect 179230 40060 179236 40072
rect 179288 40060 179294 40112
rect 182174 40060 182180 40112
rect 182232 40100 182238 40112
rect 183370 40100 183376 40112
rect 182232 40072 183376 40100
rect 182232 40060 182238 40072
rect 183370 40060 183376 40072
rect 183428 40060 183434 40112
rect 189166 40060 189172 40112
rect 189224 40100 189230 40112
rect 190362 40100 190368 40112
rect 189224 40072 190368 40100
rect 189224 40060 189230 40072
rect 190362 40060 190368 40072
rect 190420 40060 190426 40112
rect 195974 40060 195980 40112
rect 196032 40100 196038 40112
rect 197170 40100 197176 40112
rect 196032 40072 197176 40100
rect 196032 40060 196038 40072
rect 197170 40060 197176 40072
rect 197228 40060 197234 40112
rect 202966 40060 202972 40112
rect 203024 40100 203030 40112
rect 204070 40100 204076 40112
rect 203024 40072 204076 40100
rect 203024 40060 203030 40072
rect 204070 40060 204076 40072
rect 204128 40060 204134 40112
rect 209774 40060 209780 40112
rect 209832 40100 209838 40112
rect 210970 40100 210976 40112
rect 209832 40072 210976 40100
rect 209832 40060 209838 40072
rect 210970 40060 210976 40072
rect 211028 40060 211034 40112
rect 212902 40060 212908 40112
rect 212960 40100 212966 40112
rect 213730 40100 213736 40112
rect 212960 40072 213736 40100
rect 212960 40060 212966 40072
rect 213730 40060 213736 40072
rect 213788 40060 213794 40112
rect 215846 40060 215852 40112
rect 215904 40100 215910 40112
rect 216582 40100 216588 40112
rect 215904 40072 216588 40100
rect 215904 40060 215910 40072
rect 216582 40060 216588 40072
rect 216640 40060 216646 40112
rect 220814 40060 220820 40112
rect 220872 40100 220878 40112
rect 222102 40100 222108 40112
rect 220872 40072 222108 40100
rect 220872 40060 220878 40072
rect 222102 40060 222108 40072
rect 222160 40060 222166 40112
rect 230566 40060 230572 40112
rect 230624 40100 230630 40112
rect 231762 40100 231768 40112
rect 230624 40072 231768 40100
rect 230624 40060 230630 40072
rect 231762 40060 231768 40072
rect 231820 40060 231826 40112
rect 243446 40060 243452 40112
rect 243504 40100 243510 40112
rect 244182 40100 244188 40112
rect 243504 40072 244188 40100
rect 243504 40060 243510 40072
rect 244182 40060 244188 40072
rect 244240 40060 244246 40112
rect 244550 40060 244556 40112
rect 244608 40100 244614 40112
rect 245470 40100 245476 40112
rect 244608 40072 245476 40100
rect 244608 40060 244614 40072
rect 245470 40060 245476 40072
rect 245528 40060 245534 40112
rect 254302 40060 254308 40112
rect 254360 40100 254366 40112
rect 255222 40100 255228 40112
rect 254360 40072 255228 40100
rect 254360 40060 254366 40072
rect 255222 40060 255228 40072
rect 255280 40060 255286 40112
rect 269206 40060 269212 40112
rect 269264 40100 269270 40112
rect 270402 40100 270408 40112
rect 269264 40072 270408 40100
rect 269264 40060 269270 40072
rect 270402 40060 270408 40072
rect 270460 40060 270466 40112
rect 279142 40060 279148 40112
rect 279200 40100 279206 40112
rect 280062 40100 280068 40112
rect 279200 40072 280068 40100
rect 279200 40060 279206 40072
rect 280062 40060 280068 40072
rect 280120 40060 280126 40112
rect 95142 39992 95148 40044
rect 95200 40032 95206 40044
rect 533338 40032 533344 40044
rect 95200 40004 533344 40032
rect 95200 39992 95206 40004
rect 533338 39992 533344 40004
rect 533396 39992 533402 40044
rect 14458 39924 14464 39976
rect 14516 39964 14522 39976
rect 264238 39964 264244 39976
rect 14516 39936 264244 39964
rect 14516 39924 14522 39936
rect 264238 39924 264244 39936
rect 264296 39924 264302 39976
rect 265158 39924 265164 39976
rect 265216 39964 265222 39976
rect 329098 39964 329104 39976
rect 265216 39936 329104 39964
rect 265216 39924 265222 39936
rect 329098 39924 329104 39936
rect 329156 39924 329162 39976
rect 81342 39856 81348 39908
rect 81400 39896 81406 39908
rect 299750 39896 299756 39908
rect 81400 39868 299756 39896
rect 81400 39856 81406 39868
rect 299750 39856 299756 39868
rect 299808 39856 299814 39908
rect 82262 39788 82268 39840
rect 82320 39828 82326 39840
rect 295978 39828 295984 39840
rect 82320 39800 295984 39828
rect 82320 39788 82326 39800
rect 295978 39788 295984 39800
rect 296036 39788 296042 39840
rect 74350 39720 74356 39772
rect 74408 39760 74414 39772
rect 284938 39760 284944 39772
rect 74408 39732 284944 39760
rect 74408 39720 74414 39732
rect 284938 39720 284944 39732
rect 284996 39720 285002 39772
rect 219710 39652 219716 39704
rect 219768 39692 219774 39704
rect 291838 39692 291844 39704
rect 219768 39664 291844 39692
rect 219768 39652 219774 39664
rect 291838 39652 291844 39664
rect 291896 39652 291902 39704
rect 60918 39380 60924 39432
rect 60976 39420 60982 39432
rect 186314 39420 186320 39432
rect 60976 39392 186320 39420
rect 60976 39380 60982 39392
rect 186314 39380 186320 39392
rect 186372 39380 186378 39432
rect 263502 39380 263508 39432
rect 263560 39420 263566 39432
rect 281994 39420 282000 39432
rect 263560 39392 282000 39420
rect 263560 39380 263566 39392
rect 281994 39380 282000 39392
rect 282052 39380 282058 39432
rect 59722 39312 59728 39364
rect 59780 39352 59786 39364
rect 390646 39352 390652 39364
rect 59780 39324 390652 39352
rect 59780 39312 59786 39324
rect 390646 39312 390652 39324
rect 390704 39312 390710 39364
rect 135073 38675 135131 38681
rect 135073 38641 135085 38675
rect 135119 38672 135131 38675
rect 135162 38672 135168 38684
rect 135119 38644 135168 38672
rect 135119 38641 135131 38644
rect 135073 38635 135131 38641
rect 135162 38632 135168 38644
rect 135220 38632 135226 38684
rect 137002 38604 137008 38616
rect 136963 38576 137008 38604
rect 137002 38564 137008 38576
rect 137060 38564 137066 38616
rect 135073 38539 135131 38545
rect 135073 38505 135085 38539
rect 135119 38536 135131 38539
rect 135162 38536 135168 38548
rect 135119 38508 135168 38536
rect 135119 38505 135131 38508
rect 135073 38499 135131 38505
rect 135162 38496 135168 38508
rect 135220 38496 135226 38548
rect 283190 38196 283196 38208
rect 278424 38168 283196 38196
rect 245562 38088 245568 38140
rect 245620 38128 245626 38140
rect 278424 38128 278452 38168
rect 283190 38156 283196 38168
rect 283248 38156 283254 38208
rect 281534 38128 281540 38140
rect 245620 38100 278452 38128
rect 278516 38100 281540 38128
rect 245620 38088 245626 38100
rect 241422 38020 241428 38072
rect 241480 38060 241486 38072
rect 278516 38060 278544 38100
rect 281534 38088 281540 38100
rect 281592 38088 281598 38140
rect 281074 38060 281080 38072
rect 241480 38032 278544 38060
rect 278608 38032 281080 38060
rect 241480 38020 241486 38032
rect 61378 37952 61384 38004
rect 61436 37992 61442 38004
rect 193214 37992 193220 38004
rect 61436 37964 193220 37992
rect 61436 37952 61442 37964
rect 193214 37952 193220 37964
rect 193272 37952 193278 38004
rect 202782 37952 202788 38004
rect 202840 37992 202846 38004
rect 278608 37992 278636 38032
rect 281074 38020 281080 38032
rect 281132 38020 281138 38072
rect 202840 37964 278636 37992
rect 202840 37952 202846 37964
rect 280982 37952 280988 38004
rect 281040 37992 281046 38004
rect 339494 37992 339500 38004
rect 281040 37964 339500 37992
rect 281040 37952 281046 37964
rect 339494 37952 339500 37964
rect 339552 37952 339558 38004
rect 59630 37884 59636 37936
rect 59688 37924 59694 37936
rect 425146 37924 425152 37936
rect 59688 37896 425152 37924
rect 59688 37884 59694 37896
rect 425146 37884 425152 37896
rect 425204 37884 425210 37936
rect 99006 37272 99012 37324
rect 99064 37312 99070 37324
rect 99282 37312 99288 37324
rect 99064 37284 99288 37312
rect 99064 37272 99070 37284
rect 99282 37272 99288 37284
rect 99340 37272 99346 37324
rect 149054 37312 149060 37324
rect 149015 37284 149060 37312
rect 149054 37272 149060 37284
rect 149112 37272 149118 37324
rect 179322 36660 179328 36712
rect 179380 36700 179386 36712
rect 281442 36700 281448 36712
rect 179380 36672 281448 36700
rect 179380 36660 179386 36672
rect 281442 36660 281448 36672
rect 281500 36660 281506 36712
rect 58434 36592 58440 36644
rect 58492 36632 58498 36644
rect 281534 36632 281540 36644
rect 58492 36604 281540 36632
rect 58492 36592 58498 36604
rect 281534 36592 281540 36604
rect 281592 36592 281598 36644
rect 60090 36524 60096 36576
rect 60148 36564 60154 36576
rect 379514 36564 379520 36576
rect 60148 36536 379520 36564
rect 60148 36524 60154 36536
rect 379514 36524 379520 36536
rect 379572 36524 379578 36576
rect 280890 36456 280896 36508
rect 280948 36496 280954 36508
rect 281350 36496 281356 36508
rect 280948 36468 281356 36496
rect 280948 36456 280954 36468
rect 281350 36456 281356 36468
rect 281408 36456 281414 36508
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 286502 35884 286508 35896
rect 3476 35856 286508 35884
rect 3476 35844 3482 35856
rect 286502 35844 286508 35856
rect 286560 35844 286566 35896
rect 58802 35300 58808 35352
rect 58860 35340 58866 35352
rect 252554 35340 252560 35352
rect 58860 35312 252560 35340
rect 58860 35300 58866 35312
rect 252554 35300 252560 35312
rect 252612 35300 252618 35352
rect 263410 35300 263416 35352
rect 263468 35340 263474 35352
rect 283742 35340 283748 35352
rect 263468 35312 283748 35340
rect 263468 35300 263474 35312
rect 283742 35300 283748 35312
rect 283800 35300 283806 35352
rect 58894 35232 58900 35284
rect 58952 35272 58958 35284
rect 340874 35272 340880 35284
rect 58952 35244 340880 35272
rect 58952 35232 58958 35244
rect 340874 35232 340880 35244
rect 340932 35232 340938 35284
rect 62298 35164 62304 35216
rect 62356 35204 62362 35216
rect 346394 35204 346400 35216
rect 62356 35176 346400 35204
rect 62356 35164 62362 35176
rect 346394 35164 346400 35176
rect 346452 35164 346458 35216
rect 62390 35096 62396 35148
rect 62448 35096 62454 35148
rect 62408 34944 62436 35096
rect 62390 34892 62396 34944
rect 62448 34892 62454 34944
rect 219342 33872 219348 33924
rect 219400 33912 219406 33924
rect 282362 33912 282368 33924
rect 219400 33884 282368 33912
rect 219400 33872 219406 33884
rect 282362 33872 282368 33884
rect 282420 33872 282426 33924
rect 59906 33804 59912 33856
rect 59964 33844 59970 33856
rect 448514 33844 448520 33856
rect 59964 33816 448520 33844
rect 59964 33804 59970 33816
rect 448514 33804 448520 33816
rect 448572 33804 448578 33856
rect 146570 33776 146576 33788
rect 146531 33748 146576 33776
rect 146570 33736 146576 33748
rect 146628 33736 146634 33788
rect 172330 33736 172336 33788
rect 172388 33776 172394 33788
rect 572714 33776 572720 33788
rect 172388 33748 572720 33776
rect 172388 33736 172394 33748
rect 572714 33736 572720 33748
rect 572772 33736 572778 33788
rect 164142 33124 164148 33176
rect 164200 33164 164206 33176
rect 168374 33164 168380 33176
rect 164200 33136 168380 33164
rect 164200 33124 164206 33136
rect 168374 33124 168380 33136
rect 168432 33124 168438 33176
rect 179138 32512 179144 32564
rect 179196 32552 179202 32564
rect 270494 32552 270500 32564
rect 179196 32524 270500 32552
rect 179196 32512 179202 32524
rect 270494 32512 270500 32524
rect 270552 32512 270558 32564
rect 64782 32444 64788 32496
rect 64840 32484 64846 32496
rect 223206 32484 223212 32496
rect 64840 32456 223212 32484
rect 64840 32444 64846 32456
rect 223206 32444 223212 32456
rect 223264 32444 223270 32496
rect 269022 32444 269028 32496
rect 269080 32484 269086 32496
rect 280890 32484 280896 32496
rect 269080 32456 280896 32484
rect 269080 32444 269086 32456
rect 280890 32444 280896 32456
rect 280948 32444 280954 32496
rect 213730 32376 213736 32428
rect 213788 32416 213794 32428
rect 483014 32416 483020 32428
rect 213788 32388 483020 32416
rect 213788 32376 213794 32388
rect 483014 32376 483020 32388
rect 483072 32376 483078 32428
rect 237650 31832 237656 31884
rect 237708 31832 237714 31884
rect 237668 31748 237696 31832
rect 237650 31696 237656 31748
rect 237708 31696 237714 31748
rect 280062 31288 280068 31340
rect 280120 31328 280126 31340
rect 287238 31328 287244 31340
rect 280120 31300 287244 31328
rect 280120 31288 280126 31300
rect 287238 31288 287244 31300
rect 287296 31288 287302 31340
rect 119890 31220 119896 31272
rect 119948 31260 119954 31272
rect 307754 31260 307760 31272
rect 119948 31232 307760 31260
rect 119948 31220 119954 31232
rect 307754 31220 307760 31232
rect 307812 31220 307818 31272
rect 58526 31152 58532 31204
rect 58584 31192 58590 31204
rect 295334 31192 295340 31204
rect 58584 31164 295340 31192
rect 58584 31152 58590 31164
rect 295334 31152 295340 31164
rect 295392 31152 295398 31204
rect 146202 31084 146208 31136
rect 146260 31124 146266 31136
rect 226334 31124 226340 31136
rect 146260 31096 226340 31124
rect 146260 31084 146266 31096
rect 226334 31084 226340 31096
rect 226392 31084 226398 31136
rect 271782 31084 271788 31136
rect 271840 31124 271846 31136
rect 546494 31124 546500 31136
rect 271840 31096 546500 31124
rect 271840 31084 271846 31096
rect 546494 31084 546500 31096
rect 546552 31084 546558 31136
rect 59078 31016 59084 31068
rect 59136 31056 59142 31068
rect 438854 31056 438860 31068
rect 59136 31028 438860 31056
rect 59136 31016 59142 31028
rect 438854 31016 438860 31028
rect 438912 31016 438918 31068
rect 223206 30268 223212 30320
rect 223264 30308 223270 30320
rect 580166 30308 580172 30320
rect 223264 30280 580172 30308
rect 223264 30268 223270 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 128262 29656 128268 29708
rect 128320 29696 128326 29708
rect 276014 29696 276020 29708
rect 128320 29668 276020 29696
rect 128320 29656 128326 29668
rect 276014 29656 276020 29668
rect 276072 29656 276078 29708
rect 268930 29588 268936 29640
rect 268988 29628 268994 29640
rect 563054 29628 563060 29640
rect 268988 29600 563060 29628
rect 268988 29588 268994 29600
rect 563054 29588 563060 29600
rect 563112 29588 563118 29640
rect 135073 29019 135131 29025
rect 135073 28985 135085 29019
rect 135119 29016 135131 29019
rect 135162 29016 135168 29028
rect 135119 28988 135168 29016
rect 135119 28985 135131 28988
rect 135073 28979 135131 28985
rect 135162 28976 135168 28988
rect 135220 28976 135226 29028
rect 137005 29019 137063 29025
rect 137005 28985 137017 29019
rect 137051 29016 137063 29019
rect 137094 29016 137100 29028
rect 137051 28988 137100 29016
rect 137051 28985 137063 28988
rect 137005 28979 137063 28985
rect 137094 28976 137100 28988
rect 137152 28976 137158 29028
rect 146573 29019 146631 29025
rect 146573 28985 146585 29019
rect 146619 29016 146631 29019
rect 146662 29016 146668 29028
rect 146619 28988 146668 29016
rect 146619 28985 146631 28988
rect 146573 28979 146631 28985
rect 146662 28976 146668 28988
rect 146720 28976 146726 29028
rect 231762 28568 231768 28620
rect 231820 28608 231826 28620
rect 313366 28608 313372 28620
rect 231820 28580 313372 28608
rect 231820 28568 231826 28580
rect 313366 28568 313372 28580
rect 313424 28568 313430 28620
rect 124122 28500 124128 28552
rect 124180 28540 124186 28552
rect 234614 28540 234620 28552
rect 124180 28512 234620 28540
rect 124180 28500 124186 28512
rect 234614 28500 234620 28512
rect 234672 28500 234678 28552
rect 153010 28432 153016 28484
rect 153068 28472 153074 28484
rect 264974 28472 264980 28484
rect 153068 28444 264980 28472
rect 153068 28432 153074 28444
rect 264974 28432 264980 28444
rect 265032 28432 265038 28484
rect 60550 28364 60556 28416
rect 60608 28404 60614 28416
rect 350534 28404 350540 28416
rect 60608 28376 350540 28404
rect 60608 28364 60614 28376
rect 350534 28364 350540 28376
rect 350592 28364 350598 28416
rect 141970 28296 141976 28348
rect 142028 28336 142034 28348
rect 484394 28336 484400 28348
rect 142028 28308 484400 28336
rect 142028 28296 142034 28308
rect 484394 28296 484400 28308
rect 484452 28296 484458 28348
rect 158530 28228 158536 28280
rect 158588 28268 158594 28280
rect 502426 28268 502432 28280
rect 158588 28240 502432 28268
rect 158588 28228 158594 28240
rect 502426 28228 502432 28240
rect 502484 28228 502490 28280
rect 99193 27591 99251 27597
rect 99193 27557 99205 27591
rect 99239 27588 99251 27591
rect 99282 27588 99288 27600
rect 99239 27560 99288 27588
rect 99239 27557 99251 27560
rect 99193 27551 99251 27557
rect 99282 27548 99288 27560
rect 99340 27548 99346 27600
rect 149054 27588 149060 27600
rect 149015 27560 149060 27588
rect 149054 27548 149060 27560
rect 149112 27548 149118 27600
rect 150618 27548 150624 27600
rect 150676 27588 150682 27600
rect 150713 27591 150771 27597
rect 150713 27588 150725 27591
rect 150676 27560 150725 27588
rect 150676 27548 150682 27560
rect 150713 27557 150725 27560
rect 150759 27557 150771 27591
rect 150713 27551 150771 27557
rect 242158 27004 242164 27056
rect 242216 27044 242222 27056
rect 283926 27044 283932 27056
rect 242216 27016 283932 27044
rect 242216 27004 242222 27016
rect 283926 27004 283932 27016
rect 283984 27004 283990 27056
rect 58710 26936 58716 26988
rect 58768 26976 58774 26988
rect 245746 26976 245752 26988
rect 58768 26948 245752 26976
rect 58768 26936 58774 26948
rect 245746 26936 245752 26948
rect 245804 26936 245810 26988
rect 70302 26868 70308 26920
rect 70360 26908 70366 26920
rect 558914 26908 558920 26920
rect 70360 26880 558920 26908
rect 70360 26868 70366 26880
rect 558914 26868 558920 26880
rect 558972 26868 558978 26920
rect 170950 25712 170956 25764
rect 171008 25752 171014 25764
rect 282086 25752 282092 25764
rect 171008 25724 282092 25752
rect 171008 25712 171014 25724
rect 282086 25712 282092 25724
rect 282144 25712 282150 25764
rect 148962 25644 148968 25696
rect 149020 25684 149026 25696
rect 281166 25684 281172 25696
rect 149020 25656 281172 25684
rect 149020 25644 149026 25656
rect 281166 25644 281172 25656
rect 281224 25644 281230 25696
rect 61194 25576 61200 25628
rect 61252 25616 61258 25628
rect 235994 25616 236000 25628
rect 61252 25588 236000 25616
rect 61252 25576 61258 25588
rect 235994 25576 236000 25588
rect 236052 25576 236058 25628
rect 241238 25576 241244 25628
rect 241296 25616 241302 25628
rect 500954 25616 500960 25628
rect 241296 25588 500960 25616
rect 241296 25576 241302 25588
rect 500954 25576 500960 25588
rect 501012 25576 501018 25628
rect 126790 25508 126796 25560
rect 126848 25548 126854 25560
rect 391934 25548 391940 25560
rect 126848 25520 391940 25548
rect 126848 25508 126854 25520
rect 391934 25508 391940 25520
rect 391992 25508 391998 25560
rect 220722 24420 220728 24472
rect 220780 24460 220786 24472
rect 283006 24460 283012 24472
rect 220780 24432 283012 24460
rect 220780 24420 220786 24432
rect 283006 24420 283012 24432
rect 283064 24420 283070 24472
rect 85482 24352 85488 24404
rect 85540 24392 85546 24404
rect 233234 24392 233240 24404
rect 85540 24364 233240 24392
rect 85540 24352 85546 24364
rect 233234 24352 233240 24364
rect 233292 24352 233298 24404
rect 148870 24284 148876 24336
rect 148928 24324 148934 24336
rect 318794 24324 318800 24336
rect 148928 24296 318800 24324
rect 148928 24284 148934 24296
rect 318794 24284 318800 24296
rect 318852 24284 318858 24336
rect 215202 24216 215208 24268
rect 215260 24256 215266 24268
rect 401594 24256 401600 24268
rect 215260 24228 401600 24256
rect 215260 24216 215266 24228
rect 401594 24216 401600 24228
rect 401652 24216 401658 24268
rect 59170 24148 59176 24200
rect 59228 24188 59234 24200
rect 280154 24188 280160 24200
rect 59228 24160 280160 24188
rect 59228 24148 59234 24160
rect 280154 24148 280160 24160
rect 280212 24148 280218 24200
rect 135070 24080 135076 24132
rect 135128 24120 135134 24132
rect 467926 24120 467932 24132
rect 135128 24092 467932 24120
rect 135128 24080 135134 24092
rect 467926 24080 467932 24092
rect 467984 24080 467990 24132
rect 176562 22992 176568 23044
rect 176620 23032 176626 23044
rect 283466 23032 283472 23044
rect 176620 23004 283472 23032
rect 176620 22992 176626 23004
rect 283466 22992 283472 23004
rect 283524 22992 283530 23044
rect 68922 22924 68928 22976
rect 68980 22964 68986 22976
rect 248414 22964 248420 22976
rect 68980 22936 248420 22964
rect 68980 22924 68986 22936
rect 248414 22924 248420 22936
rect 248472 22924 248478 22976
rect 130930 22856 130936 22908
rect 130988 22896 130994 22908
rect 336734 22896 336740 22908
rect 130988 22868 336740 22896
rect 130988 22856 130994 22868
rect 336734 22856 336740 22868
rect 336792 22856 336798 22908
rect 60826 22788 60832 22840
rect 60884 22828 60890 22840
rect 324314 22828 324320 22840
rect 60884 22800 324320 22828
rect 60884 22788 60890 22800
rect 324314 22788 324320 22800
rect 324372 22788 324378 22840
rect 144822 22720 144828 22772
rect 144880 22760 144886 22772
rect 466454 22760 466460 22772
rect 144880 22732 466460 22760
rect 144880 22720 144886 22732
rect 466454 22720 466460 22732
rect 466512 22720 466518 22772
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 146662 22080 146668 22092
rect 3200 22052 146668 22080
rect 3200 22040 3206 22052
rect 146662 22040 146668 22052
rect 146720 22040 146726 22092
rect 139210 21496 139216 21548
rect 139268 21536 139274 21548
rect 252646 21536 252652 21548
rect 139268 21508 252652 21536
rect 139268 21496 139274 21508
rect 252646 21496 252652 21508
rect 252704 21496 252710 21548
rect 253842 21496 253848 21548
rect 253900 21536 253906 21548
rect 320174 21536 320180 21548
rect 253900 21508 320180 21536
rect 253900 21496 253906 21508
rect 320174 21496 320180 21508
rect 320232 21496 320238 21548
rect 162670 21428 162676 21480
rect 162728 21468 162734 21480
rect 282270 21468 282276 21480
rect 162728 21440 282276 21468
rect 162728 21428 162734 21440
rect 282270 21428 282276 21440
rect 282328 21428 282334 21480
rect 131022 21360 131028 21412
rect 131080 21400 131086 21412
rect 546586 21400 546592 21412
rect 131080 21372 546592 21400
rect 131080 21360 131086 21372
rect 546586 21360 546592 21372
rect 546644 21360 546650 21412
rect 203978 20000 203984 20052
rect 204036 20040 204042 20052
rect 280614 20040 280620 20052
rect 204036 20012 280620 20040
rect 204036 20000 204042 20012
rect 280614 20000 280620 20012
rect 280672 20000 280678 20052
rect 62390 19932 62396 19984
rect 62448 19972 62454 19984
rect 162854 19972 162860 19984
rect 62448 19944 162860 19972
rect 62448 19932 62454 19944
rect 162854 19932 162860 19944
rect 162912 19932 162918 19984
rect 179230 19932 179236 19984
rect 179288 19972 179294 19984
rect 516134 19972 516140 19984
rect 179288 19944 516140 19972
rect 179288 19932 179294 19944
rect 516134 19932 516140 19944
rect 516192 19932 516198 19984
rect 135162 19592 135168 19644
rect 135220 19592 135226 19644
rect 135180 19372 135208 19592
rect 135162 19320 135168 19372
rect 135220 19320 135226 19372
rect 135162 19224 135168 19236
rect 135123 19196 135168 19224
rect 135162 19184 135168 19196
rect 135220 19184 135226 19236
rect 129642 18844 129648 18896
rect 129700 18884 129706 18896
rect 237558 18884 237564 18896
rect 129700 18856 237564 18884
rect 129700 18844 129706 18856
rect 237558 18844 237564 18856
rect 237616 18844 237622 18896
rect 143350 18776 143356 18828
rect 143408 18816 143414 18828
rect 281626 18816 281632 18828
rect 143408 18788 281632 18816
rect 143408 18776 143414 18788
rect 281626 18776 281632 18788
rect 281684 18776 281690 18828
rect 182082 18708 182088 18760
rect 182140 18748 182146 18760
rect 520366 18748 520372 18760
rect 182140 18720 520372 18748
rect 182140 18708 182146 18720
rect 520366 18708 520372 18720
rect 520424 18708 520430 18760
rect 175182 18640 175188 18692
rect 175240 18680 175246 18692
rect 514754 18680 514760 18692
rect 175240 18652 514760 18680
rect 175240 18640 175246 18652
rect 514754 18640 514760 18652
rect 514812 18640 514818 18692
rect 58986 18572 58992 18624
rect 59044 18612 59050 18624
rect 488534 18612 488540 18624
rect 59044 18584 488540 18612
rect 59044 18572 59050 18584
rect 488534 18572 488540 18584
rect 488592 18572 488598 18624
rect 149054 18000 149060 18012
rect 149015 17972 149060 18000
rect 149054 17960 149060 17972
rect 149112 17960 149118 18012
rect 55950 17892 55956 17944
rect 56008 17932 56014 17944
rect 579798 17932 579804 17944
rect 56008 17904 579804 17932
rect 56008 17892 56014 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 168190 17484 168196 17536
rect 168248 17524 168254 17536
rect 269114 17524 269120 17536
rect 168248 17496 269120 17524
rect 168248 17484 168254 17496
rect 269114 17484 269120 17496
rect 269172 17484 269178 17536
rect 204070 17416 204076 17468
rect 204128 17456 204134 17468
rect 532694 17456 532700 17468
rect 204128 17428 532700 17456
rect 204128 17416 204134 17428
rect 532694 17416 532700 17428
rect 532752 17416 532758 17468
rect 57514 17348 57520 17400
rect 57572 17388 57578 17400
rect 443086 17388 443092 17400
rect 57572 17360 443092 17388
rect 57572 17348 57578 17360
rect 443086 17348 443092 17360
rect 443144 17348 443150 17400
rect 111702 17280 111708 17332
rect 111760 17320 111766 17332
rect 505094 17320 505100 17332
rect 111760 17292 505100 17320
rect 111760 17280 111766 17292
rect 505094 17280 505100 17292
rect 505152 17280 505158 17332
rect 103422 17212 103428 17264
rect 103480 17252 103486 17264
rect 513374 17252 513380 17264
rect 103480 17224 513380 17252
rect 103480 17212 103486 17224
rect 513374 17212 513380 17224
rect 513432 17212 513438 17264
rect 231762 16124 231768 16176
rect 231820 16164 231826 16176
rect 283558 16164 283564 16176
rect 231820 16136 283564 16164
rect 231820 16124 231826 16136
rect 283558 16124 283564 16136
rect 283616 16124 283622 16176
rect 118602 16056 118608 16108
rect 118660 16096 118666 16108
rect 247126 16096 247132 16108
rect 118660 16068 247132 16096
rect 118660 16056 118666 16068
rect 247126 16056 247132 16068
rect 247184 16056 247190 16108
rect 270402 16056 270408 16108
rect 270460 16096 270466 16108
rect 291194 16096 291200 16108
rect 270460 16068 291200 16096
rect 270460 16056 270466 16068
rect 291194 16056 291200 16068
rect 291252 16056 291258 16108
rect 304258 16056 304264 16108
rect 304316 16096 304322 16108
rect 528646 16096 528652 16108
rect 304316 16068 528652 16096
rect 304316 16056 304322 16068
rect 528646 16056 528652 16068
rect 528704 16056 528710 16108
rect 59262 15988 59268 16040
rect 59320 16028 59326 16040
rect 309134 16028 309140 16040
rect 59320 16000 309140 16028
rect 59320 15988 59326 16000
rect 309134 15988 309140 16000
rect 309192 15988 309198 16040
rect 115842 15920 115848 15972
rect 115900 15960 115906 15972
rect 414014 15960 414020 15972
rect 115900 15932 414020 15960
rect 115900 15920 115906 15932
rect 414014 15920 414020 15932
rect 414072 15920 414078 15972
rect 197170 15852 197176 15904
rect 197228 15892 197234 15904
rect 510614 15892 510620 15904
rect 197228 15864 510620 15892
rect 197228 15852 197234 15864
rect 510614 15852 510620 15864
rect 510672 15852 510678 15904
rect 210970 14628 210976 14680
rect 211028 14668 211034 14680
rect 321554 14668 321560 14680
rect 211028 14640 321560 14668
rect 211028 14628 211034 14640
rect 321554 14628 321560 14640
rect 321612 14628 321618 14680
rect 71590 14560 71596 14612
rect 71648 14600 71654 14612
rect 236086 14600 236092 14612
rect 71648 14572 236092 14600
rect 71648 14560 71654 14572
rect 236086 14560 236092 14572
rect 236144 14560 236150 14612
rect 240042 14560 240048 14612
rect 240100 14600 240106 14612
rect 281258 14600 281264 14612
rect 240100 14572 281264 14600
rect 240100 14560 240106 14572
rect 281258 14560 281264 14572
rect 281316 14560 281322 14612
rect 140682 14492 140688 14544
rect 140740 14532 140746 14544
rect 371234 14532 371240 14544
rect 140740 14504 371240 14532
rect 140740 14492 140746 14504
rect 371234 14492 371240 14504
rect 371292 14492 371298 14544
rect 121362 14424 121368 14476
rect 121420 14464 121426 14476
rect 569954 14464 569960 14476
rect 121420 14436 569960 14464
rect 121420 14424 121426 14436
rect 569954 14424 569960 14436
rect 570012 14424 570018 14476
rect 182082 13744 182088 13796
rect 182140 13784 182146 13796
rect 185118 13784 185124 13796
rect 182140 13756 185124 13784
rect 182140 13744 182146 13756
rect 185118 13744 185124 13756
rect 185176 13744 185182 13796
rect 256510 13200 256516 13252
rect 256568 13240 256574 13252
rect 283374 13240 283380 13252
rect 256568 13212 283380 13240
rect 256568 13200 256574 13212
rect 283374 13200 283380 13212
rect 283432 13200 283438 13252
rect 190362 13132 190368 13184
rect 190420 13172 190426 13184
rect 343634 13172 343640 13184
rect 190420 13144 343640 13172
rect 190420 13132 190426 13144
rect 343634 13132 343640 13144
rect 343692 13132 343698 13184
rect 137922 13064 137928 13116
rect 137980 13104 137986 13116
rect 553394 13104 553400 13116
rect 137980 13076 553400 13104
rect 137980 13064 137986 13076
rect 553394 13064 553400 13076
rect 553452 13064 553458 13116
rect 554038 13064 554044 13116
rect 554096 13104 554102 13116
rect 560294 13104 560300 13116
rect 554096 13076 560300 13104
rect 554096 13064 554102 13076
rect 560294 13064 560300 13076
rect 560352 13064 560358 13116
rect 149054 12452 149060 12504
rect 149112 12452 149118 12504
rect 237466 12452 237472 12504
rect 237524 12492 237530 12504
rect 237742 12492 237748 12504
rect 237524 12464 237748 12492
rect 237524 12452 237530 12464
rect 237742 12452 237748 12464
rect 237800 12452 237806 12504
rect 149072 12288 149100 12452
rect 149238 12288 149244 12300
rect 149072 12260 149244 12288
rect 149238 12248 149244 12260
rect 149296 12248 149302 12300
rect 166902 12044 166908 12096
rect 166960 12084 166966 12096
rect 247034 12084 247040 12096
rect 166960 12056 247040 12084
rect 166960 12044 166966 12056
rect 247034 12044 247040 12056
rect 247092 12044 247098 12096
rect 136450 11976 136456 12028
rect 136508 12016 136514 12028
rect 166994 12016 167000 12028
rect 136508 11988 167000 12016
rect 136508 11976 136514 11988
rect 166994 11976 167000 11988
rect 167052 11976 167058 12028
rect 183370 11976 183376 12028
rect 183428 12016 183434 12028
rect 283006 12016 283012 12028
rect 183428 11988 283012 12016
rect 183428 11976 183434 11988
rect 283006 11976 283012 11988
rect 283064 11976 283070 12028
rect 131390 11908 131396 11960
rect 131448 11948 131454 11960
rect 281902 11948 281908 11960
rect 131448 11920 281908 11948
rect 131448 11908 131454 11920
rect 281902 11908 281908 11920
rect 281960 11908 281966 11960
rect 133598 11840 133604 11892
rect 133656 11880 133662 11892
rect 237466 11880 237472 11892
rect 133656 11852 237472 11880
rect 133656 11840 133662 11852
rect 237466 11840 237472 11852
rect 237524 11840 237530 11892
rect 252462 11840 252468 11892
rect 252520 11880 252526 11892
rect 408586 11880 408592 11892
rect 252520 11852 408592 11880
rect 252520 11840 252526 11852
rect 408586 11840 408592 11852
rect 408644 11840 408650 11892
rect 60734 11772 60740 11824
rect 60792 11812 60798 11824
rect 299474 11812 299480 11824
rect 60792 11784 299480 11812
rect 60792 11772 60798 11784
rect 299474 11772 299480 11784
rect 299532 11772 299538 11824
rect 308398 11772 308404 11824
rect 308456 11812 308462 11824
rect 507854 11812 507860 11824
rect 308456 11784 507860 11812
rect 308456 11772 308462 11784
rect 507854 11772 507860 11784
rect 507912 11772 507918 11824
rect 58618 11704 58624 11756
rect 58676 11744 58682 11756
rect 444374 11744 444380 11756
rect 58676 11716 444380 11744
rect 58676 11704 58682 11716
rect 444374 11704 444380 11716
rect 444432 11704 444438 11756
rect 150710 11676 150716 11688
rect 150671 11648 150716 11676
rect 150710 11636 150716 11648
rect 150768 11636 150774 11688
rect 385678 10956 385684 11008
rect 385736 10996 385742 11008
rect 389174 10996 389180 11008
rect 385736 10968 389180 10996
rect 385736 10956 385742 10968
rect 389174 10956 389180 10968
rect 389232 10956 389238 11008
rect 409138 10956 409144 11008
rect 409196 10996 409202 11008
rect 409874 10996 409880 11008
rect 409196 10968 409880 10996
rect 409196 10956 409202 10968
rect 409874 10956 409880 10968
rect 409932 10956 409938 11008
rect 205542 10684 205548 10736
rect 205600 10724 205606 10736
rect 335354 10724 335360 10736
rect 205600 10696 335360 10724
rect 205600 10684 205606 10696
rect 335354 10684 335360 10696
rect 335412 10684 335418 10736
rect 172422 10616 172428 10668
rect 172480 10656 172486 10668
rect 342254 10656 342260 10668
rect 172480 10628 342260 10656
rect 172480 10616 172486 10628
rect 342254 10616 342260 10628
rect 342312 10616 342318 10668
rect 193122 10548 193128 10600
rect 193180 10588 193186 10600
rect 364334 10588 364340 10600
rect 193180 10560 364340 10588
rect 193180 10548 193186 10560
rect 364334 10548 364340 10560
rect 364392 10548 364398 10600
rect 171042 10480 171048 10532
rect 171100 10520 171106 10532
rect 353294 10520 353300 10532
rect 171100 10492 353300 10520
rect 171100 10480 171106 10492
rect 353294 10480 353300 10492
rect 353352 10480 353358 10532
rect 155770 10412 155776 10464
rect 155828 10452 155834 10464
rect 349154 10452 349160 10464
rect 155828 10424 349160 10452
rect 155828 10412 155834 10424
rect 349154 10412 349160 10424
rect 349212 10412 349218 10464
rect 371878 10412 371884 10464
rect 371936 10452 371942 10464
rect 385034 10452 385040 10464
rect 371936 10424 385040 10452
rect 371936 10412 371942 10424
rect 385034 10412 385040 10424
rect 385092 10412 385098 10464
rect 92290 10344 92296 10396
rect 92348 10384 92354 10396
rect 356146 10384 356152 10396
rect 92348 10356 356152 10384
rect 92348 10344 92354 10356
rect 356146 10344 356152 10356
rect 356204 10344 356210 10396
rect 364978 10344 364984 10396
rect 365036 10384 365042 10396
rect 382274 10384 382280 10396
rect 365036 10356 382280 10384
rect 365036 10344 365042 10356
rect 382274 10344 382280 10356
rect 382332 10344 382338 10396
rect 389818 10344 389824 10396
rect 389876 10384 389882 10396
rect 407114 10384 407120 10396
rect 389876 10356 407120 10384
rect 389876 10344 389882 10356
rect 407114 10344 407120 10356
rect 407172 10344 407178 10396
rect 60642 10276 60648 10328
rect 60700 10316 60706 10328
rect 328454 10316 328460 10328
rect 60700 10288 328460 10316
rect 60700 10276 60706 10288
rect 328454 10276 328460 10288
rect 328512 10276 328518 10328
rect 356698 10276 356704 10328
rect 356756 10316 356762 10328
rect 463694 10316 463700 10328
rect 356756 10288 463700 10316
rect 356756 10276 356762 10288
rect 463694 10276 463700 10288
rect 463752 10276 463758 10328
rect 99190 9704 99196 9716
rect 99151 9676 99196 9704
rect 99190 9664 99196 9676
rect 99248 9664 99254 9716
rect 134886 9664 134892 9716
rect 134944 9704 134950 9716
rect 135165 9707 135223 9713
rect 135165 9704 135177 9707
rect 134944 9676 135177 9704
rect 134944 9664 134950 9676
rect 135165 9673 135177 9676
rect 135211 9673 135223 9707
rect 135165 9667 135223 9673
rect 234522 9664 234528 9716
rect 234580 9704 234586 9716
rect 234798 9704 234804 9716
rect 234580 9676 234804 9704
rect 234580 9664 234586 9676
rect 234798 9664 234804 9676
rect 234856 9664 234862 9716
rect 169662 9596 169668 9648
rect 169720 9636 169726 9648
rect 250346 9636 250352 9648
rect 169720 9608 250352 9636
rect 169720 9596 169726 9608
rect 250346 9596 250352 9608
rect 250404 9596 250410 9648
rect 257430 9596 257436 9648
rect 257488 9636 257494 9648
rect 288618 9636 288624 9648
rect 257488 9608 288624 9636
rect 257488 9596 257494 9608
rect 288618 9596 288624 9608
rect 288676 9596 288682 9648
rect 162762 9528 162768 9580
rect 162820 9568 162826 9580
rect 243170 9568 243176 9580
rect 162820 9540 243176 9568
rect 162820 9528 162826 9540
rect 243170 9528 243176 9540
rect 243228 9528 243234 9580
rect 245470 9528 245476 9580
rect 245528 9568 245534 9580
rect 303798 9568 303804 9580
rect 245528 9540 303804 9568
rect 245528 9528 245534 9540
rect 303798 9528 303804 9540
rect 303856 9528 303862 9580
rect 187602 9460 187608 9512
rect 187660 9500 187666 9512
rect 318058 9500 318064 9512
rect 187660 9472 318064 9500
rect 187660 9460 187666 9472
rect 318058 9460 318064 9472
rect 318116 9460 318122 9512
rect 122742 9392 122748 9444
rect 122800 9432 122806 9444
rect 275278 9432 275284 9444
rect 122800 9404 275284 9432
rect 122800 9392 122806 9404
rect 275278 9392 275284 9404
rect 275336 9392 275342 9444
rect 113082 9324 113088 9376
rect 113140 9364 113146 9376
rect 321646 9364 321652 9376
rect 113140 9336 321652 9364
rect 113140 9324 113146 9336
rect 321646 9324 321652 9336
rect 321704 9324 321710 9376
rect 53374 9256 53380 9308
rect 53432 9296 53438 9308
rect 278866 9296 278872 9308
rect 53432 9268 278872 9296
rect 53432 9256 53438 9268
rect 278866 9256 278872 9268
rect 278924 9256 278930 9308
rect 180702 9188 180708 9240
rect 180760 9228 180766 9240
rect 225322 9228 225328 9240
rect 180760 9200 225328 9228
rect 180760 9188 180766 9200
rect 225322 9188 225328 9200
rect 225380 9188 225386 9240
rect 239398 9188 239404 9240
rect 239456 9228 239462 9240
rect 478690 9228 478696 9240
rect 239456 9200 478696 9228
rect 239456 9188 239462 9200
rect 478690 9188 478696 9200
rect 478748 9188 478754 9240
rect 53190 9120 53196 9172
rect 53248 9160 53254 9172
rect 294322 9160 294328 9172
rect 53248 9132 294328 9160
rect 53248 9120 53254 9132
rect 294322 9120 294328 9132
rect 294380 9120 294386 9172
rect 54662 9052 54668 9104
rect 54720 9092 54726 9104
rect 315758 9092 315764 9104
rect 54720 9064 315764 9092
rect 54720 9052 54726 9064
rect 315758 9052 315764 9064
rect 315816 9052 315822 9104
rect 322198 9052 322204 9104
rect 322256 9092 322262 9104
rect 360930 9092 360936 9104
rect 322256 9064 360936 9092
rect 322256 9052 322262 9064
rect 360930 9052 360936 9064
rect 360988 9052 360994 9104
rect 53282 8984 53288 9036
rect 53340 9024 53346 9036
rect 326430 9024 326436 9036
rect 53340 8996 326436 9024
rect 53340 8984 53346 8996
rect 326430 8984 326436 8996
rect 326488 8984 326494 9036
rect 126882 8916 126888 8968
rect 126940 8956 126946 8968
rect 228910 8956 228916 8968
rect 126940 8928 228916 8956
rect 126940 8916 126946 8928
rect 228910 8916 228916 8928
rect 228968 8916 228974 8968
rect 256602 8916 256608 8968
rect 256660 8956 256666 8968
rect 575014 8956 575020 8968
rect 256660 8928 575020 8956
rect 256660 8916 256666 8928
rect 575014 8916 575020 8928
rect 575072 8916 575078 8968
rect 196802 8848 196808 8900
rect 196860 8888 196866 8900
rect 251174 8888 251180 8900
rect 196860 8860 251180 8888
rect 196860 8848 196866 8860
rect 251174 8848 251180 8860
rect 251232 8848 251238 8900
rect 264606 8848 264612 8900
rect 264664 8888 264670 8900
rect 289814 8888 289820 8900
rect 264664 8860 289820 8888
rect 264664 8848 264670 8860
rect 289814 8848 289820 8860
rect 289872 8848 289878 8900
rect 189626 8780 189632 8832
rect 189684 8820 189690 8832
rect 241514 8820 241520 8832
rect 189684 8792 241520 8820
rect 189684 8780 189690 8792
rect 241514 8780 241520 8792
rect 241572 8780 241578 8832
rect 218146 8712 218152 8764
rect 218204 8752 218210 8764
rect 237374 8752 237380 8764
rect 218204 8724 237380 8752
rect 218204 8712 218210 8724
rect 237374 8712 237380 8724
rect 237432 8712 237438 8764
rect 208210 7964 208216 8016
rect 208268 8004 208274 8016
rect 214650 8004 214656 8016
rect 208268 7976 214656 8004
rect 208268 7964 208274 7976
rect 214650 7964 214656 7976
rect 214708 7964 214714 8016
rect 159910 7896 159916 7948
rect 159968 7936 159974 7948
rect 282914 7936 282920 7948
rect 159968 7908 282920 7936
rect 159968 7896 159974 7908
rect 282914 7896 282920 7908
rect 282972 7896 282978 7948
rect 184842 7828 184848 7880
rect 184900 7868 184906 7880
rect 395430 7868 395436 7880
rect 184900 7840 395436 7868
rect 184900 7828 184906 7840
rect 395430 7828 395436 7840
rect 395488 7828 395494 7880
rect 61102 7760 61108 7812
rect 61160 7800 61166 7812
rect 221734 7800 221740 7812
rect 61160 7772 221740 7800
rect 61160 7760 61166 7772
rect 221734 7760 221740 7772
rect 221792 7760 221798 7812
rect 224862 7760 224868 7812
rect 224920 7800 224926 7812
rect 545298 7800 545304 7812
rect 224920 7772 545304 7800
rect 224920 7760 224926 7772
rect 545298 7760 545304 7772
rect 545356 7760 545362 7812
rect 213822 7692 213828 7744
rect 213880 7732 213886 7744
rect 538122 7732 538128 7744
rect 213880 7704 538128 7732
rect 213880 7692 213886 7704
rect 538122 7692 538128 7704
rect 538180 7692 538186 7744
rect 65518 7624 65524 7676
rect 65576 7664 65582 7676
rect 399018 7664 399024 7676
rect 65576 7636 399024 7664
rect 65576 7624 65582 7636
rect 399018 7624 399024 7636
rect 399076 7624 399082 7676
rect 204162 7556 204168 7608
rect 204220 7596 204226 7608
rect 555970 7596 555976 7608
rect 204220 7568 555976 7596
rect 204220 7556 204226 7568
rect 555970 7556 555976 7568
rect 556028 7556 556034 7608
rect 2958 7352 2964 7404
rect 3016 7392 3022 7404
rect 6178 7392 6184 7404
rect 3016 7364 6184 7392
rect 3016 7352 3022 7364
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 212258 6808 212264 6860
rect 212316 6848 212322 6860
rect 284570 6848 284576 6860
rect 212316 6820 284576 6848
rect 212316 6808 212322 6820
rect 284570 6808 284576 6820
rect 284628 6808 284634 6860
rect 192018 6740 192024 6792
rect 192076 6780 192082 6792
rect 281810 6780 281816 6792
rect 192076 6752 281816 6780
rect 192076 6740 192082 6752
rect 281810 6740 281816 6752
rect 281868 6740 281874 6792
rect 144454 6672 144460 6724
rect 144512 6712 144518 6724
rect 223666 6712 223672 6724
rect 144512 6684 223672 6712
rect 144512 6672 144518 6684
rect 223666 6672 223672 6684
rect 223724 6672 223730 6724
rect 251082 6672 251088 6724
rect 251140 6712 251146 6724
rect 388254 6712 388260 6724
rect 251140 6684 388260 6712
rect 251140 6672 251146 6684
rect 388254 6672 388260 6684
rect 388312 6672 388318 6724
rect 53650 6604 53656 6656
rect 53708 6644 53714 6656
rect 177758 6644 177764 6656
rect 53708 6616 177764 6644
rect 53708 6604 53714 6616
rect 177758 6604 177764 6616
rect 177816 6604 177822 6656
rect 182542 6604 182548 6656
rect 182600 6644 182606 6656
rect 245654 6644 245660 6656
rect 182600 6616 245660 6644
rect 182600 6604 182606 6616
rect 245654 6604 245660 6616
rect 245712 6604 245718 6656
rect 266170 6604 266176 6656
rect 266228 6644 266234 6656
rect 404906 6644 404912 6656
rect 266228 6616 404912 6644
rect 266228 6604 266234 6616
rect 404906 6604 404912 6616
rect 404964 6604 404970 6656
rect 54846 6536 54852 6588
rect 54904 6576 54910 6588
rect 272886 6576 272892 6588
rect 54904 6548 272892 6576
rect 54904 6536 54910 6548
rect 272886 6536 272892 6548
rect 272944 6536 272950 6588
rect 274542 6536 274548 6588
rect 274600 6576 274606 6588
rect 365806 6576 365812 6588
rect 274600 6548 365812 6576
rect 274600 6536 274606 6548
rect 365806 6536 365812 6548
rect 365864 6536 365870 6588
rect 55674 6468 55680 6520
rect 55732 6508 55738 6520
rect 279970 6508 279976 6520
rect 55732 6480 279976 6508
rect 55732 6468 55738 6480
rect 279970 6468 279976 6480
rect 280028 6468 280034 6520
rect 53742 6400 53748 6452
rect 53800 6440 53806 6452
rect 195606 6440 195612 6452
rect 53800 6412 195612 6440
rect 53800 6400 53806 6412
rect 195606 6400 195612 6412
rect 195664 6400 195670 6452
rect 226242 6400 226248 6452
rect 226300 6440 226306 6452
rect 495342 6440 495348 6452
rect 226300 6412 495348 6440
rect 226300 6400 226306 6412
rect 495342 6400 495348 6412
rect 495400 6400 495406 6452
rect 133782 6332 133788 6384
rect 133840 6372 133846 6384
rect 422754 6372 422760 6384
rect 133840 6344 422760 6372
rect 133840 6332 133846 6344
rect 422754 6332 422760 6344
rect 422812 6332 422818 6384
rect 92382 6264 92388 6316
rect 92440 6304 92446 6316
rect 383562 6304 383568 6316
rect 92440 6276 383568 6304
rect 92440 6264 92446 6276
rect 383562 6264 383568 6276
rect 383620 6264 383626 6316
rect 54938 6196 54944 6248
rect 54996 6236 55002 6248
rect 213454 6236 213460 6248
rect 54996 6208 213460 6236
rect 54996 6196 55002 6208
rect 213454 6196 213460 6208
rect 213512 6196 213518 6248
rect 241330 6196 241336 6248
rect 241388 6236 241394 6248
rect 541710 6236 541716 6248
rect 241388 6208 541716 6236
rect 241388 6196 241394 6208
rect 541710 6196 541716 6208
rect 541768 6196 541774 6248
rect 119982 6128 119988 6180
rect 120040 6168 120046 6180
rect 440602 6168 440608 6180
rect 120040 6140 440608 6168
rect 120040 6128 120046 6140
rect 440602 6128 440608 6140
rect 440660 6128 440666 6180
rect 244182 6060 244188 6112
rect 244240 6100 244246 6112
rect 306190 6100 306196 6112
rect 244240 6072 306196 6100
rect 244240 6060 244246 6072
rect 306190 6060 306196 6072
rect 306248 6060 306254 6112
rect 266998 5992 267004 6044
rect 267056 6032 267062 6044
rect 284386 6032 284392 6044
rect 267056 6004 284392 6032
rect 267056 5992 267062 6004
rect 284386 5992 284392 6004
rect 284444 5992 284450 6044
rect 277670 5924 277676 5976
rect 277728 5964 277734 5976
rect 288526 5964 288532 5976
rect 277728 5936 288532 5964
rect 277728 5924 277734 5936
rect 288526 5924 288532 5936
rect 288584 5924 288590 5976
rect 180150 5176 180156 5228
rect 180208 5216 180214 5228
rect 198734 5216 198740 5228
rect 180208 5188 198740 5216
rect 180208 5176 180214 5188
rect 198734 5176 198740 5188
rect 198792 5176 198798 5228
rect 183462 5108 183468 5160
rect 183520 5148 183526 5160
rect 215846 5148 215852 5160
rect 183520 5120 215852 5148
rect 183520 5108 183526 5120
rect 215846 5108 215852 5120
rect 215904 5108 215910 5160
rect 222102 5108 222108 5160
rect 222160 5148 222166 5160
rect 230106 5148 230112 5160
rect 222160 5120 230112 5148
rect 222160 5108 222166 5120
rect 230106 5108 230112 5120
rect 230164 5108 230170 5160
rect 241974 5108 241980 5160
rect 242032 5148 242038 5160
rect 283650 5148 283656 5160
rect 242032 5120 283656 5148
rect 242032 5108 242038 5120
rect 283650 5108 283656 5120
rect 283708 5108 283714 5160
rect 132402 5040 132408 5092
rect 132460 5080 132466 5092
rect 201494 5080 201500 5092
rect 132460 5052 201500 5080
rect 132460 5040 132466 5052
rect 201494 5040 201500 5052
rect 201552 5040 201558 5092
rect 208670 5040 208676 5092
rect 208728 5080 208734 5092
rect 260834 5080 260840 5092
rect 208728 5052 260840 5080
rect 208728 5040 208734 5052
rect 260834 5040 260840 5052
rect 260892 5040 260898 5092
rect 267642 5040 267648 5092
rect 267700 5080 267706 5092
rect 271690 5080 271696 5092
rect 267700 5052 271696 5080
rect 267700 5040 267706 5052
rect 271690 5040 271696 5052
rect 271748 5040 271754 5092
rect 143442 4972 143448 5024
rect 143500 5012 143506 5024
rect 274082 5012 274088 5024
rect 143500 4984 274088 5012
rect 143500 4972 143506 4984
rect 274082 4972 274088 4984
rect 274140 4972 274146 5024
rect 278682 4972 278688 5024
rect 278740 5012 278746 5024
rect 551186 5012 551192 5024
rect 278740 4984 551192 5012
rect 278740 4972 278746 4984
rect 551186 4972 551192 4984
rect 551244 4972 551250 5024
rect 197262 4904 197268 4956
rect 197320 4944 197326 4956
rect 523862 4944 523868 4956
rect 197320 4916 523868 4944
rect 197320 4904 197326 4916
rect 523862 4904 523868 4916
rect 523920 4904 523926 4956
rect 108942 4836 108948 4888
rect 109000 4876 109006 4888
rect 453666 4876 453672 4888
rect 109000 4848 453672 4876
rect 109000 4836 109006 4848
rect 453666 4836 453672 4848
rect 453724 4836 453730 4888
rect 71682 4768 71688 4820
rect 71740 4808 71746 4820
rect 579798 4808 579804 4820
rect 71740 4780 579804 4808
rect 71740 4768 71746 4780
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 281534 4156 281540 4208
rect 281592 4196 281598 4208
rect 282454 4196 282460 4208
rect 281592 4168 282460 4196
rect 281592 4156 281598 4168
rect 282454 4156 282460 4168
rect 282512 4156 282518 4208
rect 55030 4088 55036 4140
rect 55088 4128 55094 4140
rect 161106 4128 161112 4140
rect 55088 4100 161112 4128
rect 55088 4088 55094 4100
rect 161106 4088 161112 4100
rect 161164 4088 161170 4140
rect 239582 4088 239588 4140
rect 239640 4128 239646 4140
rect 240042 4128 240048 4140
rect 239640 4100 240048 4128
rect 239640 4088 239646 4100
rect 240042 4088 240048 4100
rect 240100 4088 240106 4140
rect 255038 4088 255044 4140
rect 255096 4128 255102 4140
rect 287146 4128 287152 4140
rect 255096 4100 287152 4128
rect 255096 4088 255102 4100
rect 287146 4088 287152 4100
rect 287204 4088 287210 4140
rect 514018 4088 514024 4140
rect 514076 4128 514082 4140
rect 514570 4128 514576 4140
rect 514076 4100 514576 4128
rect 514076 4088 514082 4100
rect 514570 4088 514576 4100
rect 514628 4088 514634 4140
rect 57790 4020 57796 4072
rect 57848 4060 57854 4072
rect 164694 4060 164700 4072
rect 57848 4032 164700 4060
rect 57848 4020 57854 4032
rect 164694 4020 164700 4032
rect 164752 4020 164758 4072
rect 205082 4020 205088 4072
rect 205140 4060 205146 4072
rect 279418 4060 279424 4072
rect 205140 4032 279424 4060
rect 205140 4020 205146 4032
rect 279418 4020 279424 4032
rect 279476 4020 279482 4072
rect 281534 4020 281540 4072
rect 281592 4060 281598 4072
rect 282178 4060 282184 4072
rect 281592 4032 282184 4060
rect 281592 4020 281598 4032
rect 282178 4020 282184 4032
rect 282236 4020 282242 4072
rect 403618 4020 403624 4072
rect 403676 4060 403682 4072
rect 409785 4063 409843 4069
rect 409785 4060 409797 4063
rect 403676 4032 409797 4060
rect 403676 4020 403682 4032
rect 409785 4029 409797 4032
rect 409831 4029 409843 4063
rect 409785 4023 409843 4029
rect 56410 3952 56416 4004
rect 56468 3992 56474 4004
rect 176470 3992 176476 4004
rect 56468 3964 176476 3992
rect 56468 3952 56474 3964
rect 176470 3952 176476 3964
rect 176528 3952 176534 4004
rect 183738 3952 183744 4004
rect 183796 3992 183802 4004
rect 285766 3992 285772 4004
rect 183796 3964 285772 3992
rect 183796 3952 183802 3964
rect 285766 3952 285772 3964
rect 285824 3952 285830 4004
rect 407758 3952 407764 4004
rect 407816 3992 407822 4004
rect 435818 3992 435824 4004
rect 407816 3964 435824 3992
rect 407816 3952 407822 3964
rect 435818 3952 435824 3964
rect 435876 3952 435882 4004
rect 57882 3884 57888 3936
rect 57940 3924 57946 3936
rect 186038 3924 186044 3936
rect 57940 3896 186044 3924
rect 57940 3884 57946 3896
rect 186038 3884 186044 3896
rect 186096 3884 186102 3936
rect 199194 3884 199200 3936
rect 199252 3924 199258 3936
rect 281718 3924 281724 3936
rect 199252 3896 281724 3924
rect 199252 3884 199258 3896
rect 281718 3884 281724 3896
rect 281776 3884 281782 3936
rect 356146 3884 356152 3936
rect 356204 3924 356210 3936
rect 357342 3924 357348 3936
rect 356204 3896 357348 3924
rect 356204 3884 356210 3896
rect 357342 3884 357348 3896
rect 357400 3884 357406 3936
rect 390646 3884 390652 3936
rect 390704 3924 390710 3936
rect 391842 3924 391848 3936
rect 390704 3896 391848 3924
rect 390704 3884 390710 3896
rect 391842 3884 391848 3896
rect 391900 3884 391906 3936
rect 408494 3884 408500 3936
rect 408552 3924 408558 3936
rect 409690 3924 409696 3936
rect 408552 3896 409696 3924
rect 408552 3884 408558 3896
rect 409690 3884 409696 3896
rect 409748 3884 409754 3936
rect 409785 3927 409843 3933
rect 409785 3893 409797 3927
rect 409831 3924 409843 3927
rect 432322 3924 432328 3936
rect 409831 3896 432328 3924
rect 409831 3893 409843 3896
rect 409785 3887 409843 3893
rect 432322 3884 432328 3896
rect 432380 3884 432386 3936
rect 57146 3816 57152 3868
rect 57204 3856 57210 3868
rect 190822 3856 190828 3868
rect 57204 3828 190828 3856
rect 57204 3816 57210 3828
rect 190822 3816 190828 3828
rect 190880 3816 190886 3868
rect 217042 3816 217048 3868
rect 217100 3856 217106 3868
rect 242158 3856 242164 3868
rect 217100 3828 242164 3856
rect 217100 3816 217106 3828
rect 242158 3816 242164 3828
rect 242216 3816 242222 3868
rect 255958 3816 255964 3868
rect 256016 3856 256022 3868
rect 417970 3856 417976 3868
rect 256016 3828 417976 3856
rect 256016 3816 256022 3828
rect 417970 3816 417976 3828
rect 418028 3816 418034 3868
rect 57606 3748 57612 3800
rect 57664 3788 57670 3800
rect 222930 3788 222936 3800
rect 57664 3760 222936 3788
rect 57664 3748 57670 3760
rect 222930 3748 222936 3760
rect 222988 3748 222994 3800
rect 255222 3748 255228 3800
rect 255280 3788 255286 3800
rect 421558 3788 421564 3800
rect 255280 3760 421564 3788
rect 255280 3748 255286 3760
rect 421558 3748 421564 3760
rect 421616 3748 421622 3800
rect 53558 3680 53564 3732
rect 53616 3720 53622 3732
rect 244366 3720 244372 3732
rect 53616 3692 244372 3720
rect 53616 3680 53622 3692
rect 244366 3680 244372 3692
rect 244424 3680 244430 3732
rect 251450 3680 251456 3732
rect 251508 3720 251514 3732
rect 284478 3720 284484 3732
rect 251508 3692 284484 3720
rect 251508 3680 251514 3692
rect 284478 3680 284484 3692
rect 284536 3680 284542 3732
rect 285214 3680 285220 3732
rect 285272 3720 285278 3732
rect 475102 3720 475108 3732
rect 285272 3692 475108 3720
rect 285272 3680 285278 3692
rect 475102 3680 475108 3692
rect 475160 3680 475166 3732
rect 502978 3680 502984 3732
rect 503036 3720 503042 3732
rect 503036 3692 503760 3720
rect 503036 3680 503042 3692
rect 57698 3612 57704 3664
rect 57756 3652 57762 3664
rect 197998 3652 198004 3664
rect 57756 3624 198004 3652
rect 57756 3612 57762 3624
rect 197998 3612 198004 3624
rect 198056 3612 198062 3664
rect 204898 3612 204904 3664
rect 204956 3652 204962 3664
rect 425054 3652 425060 3664
rect 204956 3624 425060 3652
rect 204956 3612 204962 3624
rect 425054 3612 425060 3624
rect 425112 3612 425118 3664
rect 459646 3612 459652 3664
rect 459704 3652 459710 3664
rect 460842 3652 460848 3664
rect 459704 3624 460848 3652
rect 459704 3612 459710 3624
rect 460842 3612 460848 3624
rect 460900 3612 460906 3664
rect 467098 3612 467104 3664
rect 467156 3652 467162 3664
rect 497734 3652 497740 3664
rect 467156 3624 497740 3652
rect 467156 3612 467162 3624
rect 497734 3612 497740 3624
rect 497792 3612 497798 3664
rect 64138 3544 64144 3596
rect 64196 3584 64202 3596
rect 206278 3584 206284 3596
rect 64196 3556 206284 3584
rect 64196 3544 64202 3556
rect 206278 3544 206284 3556
rect 206336 3544 206342 3596
rect 216582 3544 216588 3596
rect 216640 3584 216646 3596
rect 471514 3584 471520 3596
rect 216640 3556 471520 3584
rect 216640 3544 216646 3556
rect 471514 3544 471520 3556
rect 471572 3544 471578 3596
rect 496078 3544 496084 3596
rect 496136 3584 496142 3596
rect 502334 3584 502340 3596
rect 496136 3556 502340 3584
rect 496136 3544 496142 3556
rect 502334 3544 502340 3556
rect 502392 3544 502398 3596
rect 502426 3544 502432 3596
rect 502484 3584 502490 3596
rect 503622 3584 503628 3596
rect 502484 3556 503628 3584
rect 502484 3544 502490 3556
rect 503622 3544 503628 3556
rect 503680 3544 503686 3596
rect 503732 3584 503760 3692
rect 520274 3612 520280 3664
rect 520332 3652 520338 3664
rect 521470 3652 521476 3664
rect 520332 3624 521476 3652
rect 520332 3612 520338 3624
rect 521470 3612 521476 3624
rect 521528 3612 521534 3664
rect 528646 3612 528652 3664
rect 528704 3652 528710 3664
rect 529842 3652 529848 3664
rect 528704 3624 529848 3652
rect 528704 3612 528710 3624
rect 529842 3612 529848 3624
rect 529900 3612 529906 3664
rect 552382 3584 552388 3596
rect 503732 3556 552388 3584
rect 552382 3544 552388 3556
rect 552440 3544 552446 3596
rect 563146 3544 563152 3596
rect 563204 3584 563210 3596
rect 564342 3584 564348 3596
rect 563204 3556 564348 3584
rect 563204 3544 563210 3556
rect 564342 3544 564348 3556
rect 564400 3544 564406 3596
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 89717 3519 89775 3525
rect 89717 3485 89729 3519
rect 89763 3516 89775 3519
rect 101401 3519 101459 3525
rect 101401 3516 101413 3519
rect 89763 3488 101413 3516
rect 89763 3485 89775 3488
rect 89717 3479 89775 3485
rect 101401 3485 101413 3488
rect 101447 3485 101459 3519
rect 101401 3479 101459 3485
rect 104161 3519 104219 3525
rect 104161 3485 104173 3519
rect 104207 3516 104219 3519
rect 104207 3488 113956 3516
rect 104207 3485 104219 3488
rect 104161 3479 104219 3485
rect 55122 3408 55128 3460
rect 55180 3448 55186 3460
rect 94501 3451 94559 3457
rect 94501 3448 94513 3451
rect 55180 3420 94513 3448
rect 55180 3408 55186 3420
rect 94501 3417 94513 3420
rect 94547 3417 94559 3451
rect 94501 3411 94559 3417
rect 62482 3340 62488 3392
rect 62540 3380 62546 3392
rect 89717 3383 89775 3389
rect 89717 3380 89729 3383
rect 62540 3352 89729 3380
rect 62540 3340 62546 3352
rect 89717 3349 89729 3352
rect 89763 3349 89775 3383
rect 113928 3380 113956 3488
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 425057 3519 425115 3525
rect 425057 3516 425069 3519
rect 115256 3488 425069 3516
rect 115256 3476 115262 3488
rect 425057 3485 425069 3488
rect 425103 3485 425115 3519
rect 425057 3479 425115 3485
rect 425146 3476 425152 3528
rect 425204 3516 425210 3528
rect 426342 3516 426348 3528
rect 425204 3488 426348 3516
rect 425204 3476 425210 3488
rect 426342 3476 426348 3488
rect 426400 3476 426406 3528
rect 433334 3476 433340 3528
rect 433392 3516 433398 3528
rect 434622 3516 434628 3528
rect 433392 3488 434628 3516
rect 433392 3476 433398 3488
rect 434622 3476 434628 3488
rect 434680 3476 434686 3528
rect 435358 3476 435364 3528
rect 435416 3516 435422 3528
rect 567838 3516 567844 3528
rect 435416 3488 567844 3516
rect 435416 3476 435422 3488
rect 567838 3476 567844 3488
rect 567896 3476 567902 3528
rect 574738 3476 574744 3528
rect 574796 3516 574802 3528
rect 580994 3516 581000 3528
rect 574796 3488 581000 3516
rect 574796 3476 574802 3488
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 128357 3451 128415 3457
rect 128357 3448 128369 3451
rect 122668 3420 128369 3448
rect 122668 3380 122696 3420
rect 128357 3417 128369 3420
rect 128403 3417 128415 3451
rect 128357 3411 128415 3417
rect 128446 3408 128452 3460
rect 128504 3448 128510 3460
rect 128998 3448 129004 3460
rect 128504 3420 129004 3448
rect 128504 3408 128510 3420
rect 128998 3408 129004 3420
rect 129056 3408 129062 3460
rect 136082 3408 136088 3460
rect 136140 3448 136146 3460
rect 136542 3448 136548 3460
rect 136140 3420 136548 3448
rect 136140 3408 136146 3420
rect 136542 3408 136548 3420
rect 136600 3408 136606 3460
rect 136726 3408 136732 3460
rect 136784 3448 136790 3460
rect 137278 3448 137284 3460
rect 136784 3420 137284 3448
rect 136784 3408 136790 3420
rect 137278 3408 137284 3420
rect 137336 3408 137342 3460
rect 138474 3408 138480 3460
rect 138532 3448 138538 3460
rect 139302 3448 139308 3460
rect 138532 3420 139308 3448
rect 138532 3408 138538 3420
rect 139302 3408 139308 3420
rect 139360 3408 139366 3460
rect 140866 3408 140872 3460
rect 140924 3448 140930 3460
rect 142062 3448 142068 3460
rect 140924 3420 142068 3448
rect 140924 3408 140930 3420
rect 142062 3408 142068 3420
rect 142120 3408 142126 3460
rect 144178 3408 144184 3460
rect 144236 3448 144242 3460
rect 145650 3448 145656 3460
rect 144236 3420 145656 3448
rect 144236 3408 144242 3420
rect 145650 3408 145656 3420
rect 145708 3408 145714 3460
rect 148042 3408 148048 3460
rect 148100 3448 148106 3460
rect 148962 3448 148968 3460
rect 148100 3420 148968 3448
rect 148100 3408 148106 3420
rect 148962 3408 148968 3420
rect 149020 3408 149026 3460
rect 150710 3408 150716 3460
rect 150768 3448 150774 3460
rect 151538 3448 151544 3460
rect 150768 3420 151544 3448
rect 150768 3408 150774 3420
rect 151538 3408 151544 3420
rect 151596 3408 151602 3460
rect 153930 3408 153936 3460
rect 153988 3448 153994 3460
rect 154482 3448 154488 3460
rect 153988 3420 154488 3448
rect 153988 3408 153994 3420
rect 154482 3408 154488 3420
rect 154540 3408 154546 3460
rect 155126 3408 155132 3460
rect 155184 3448 155190 3460
rect 155862 3448 155868 3460
rect 155184 3420 155868 3448
rect 155184 3408 155190 3420
rect 155862 3408 155868 3420
rect 155920 3408 155926 3460
rect 482278 3448 482284 3460
rect 155972 3420 482284 3448
rect 113928 3352 122696 3380
rect 89717 3343 89775 3349
rect 122742 3340 122748 3392
rect 122800 3380 122806 3392
rect 122800 3352 130148 3380
rect 122800 3340 122806 3352
rect 56502 3272 56508 3324
rect 56560 3312 56566 3324
rect 108945 3315 109003 3321
rect 108945 3312 108957 3315
rect 56560 3284 108957 3312
rect 56560 3272 56566 3284
rect 108945 3281 108957 3284
rect 108991 3281 109003 3315
rect 108945 3275 109003 3281
rect 109037 3315 109095 3321
rect 109037 3281 109049 3315
rect 109083 3312 109095 3315
rect 109083 3284 126560 3312
rect 109083 3281 109095 3284
rect 109037 3275 109095 3281
rect 101401 3247 101459 3253
rect 101401 3213 101413 3247
rect 101447 3244 101459 3247
rect 106277 3247 106335 3253
rect 106277 3244 106289 3247
rect 101447 3216 106289 3244
rect 101447 3213 101459 3216
rect 101401 3207 101459 3213
rect 106277 3213 106289 3216
rect 106323 3213 106335 3247
rect 106277 3207 106335 3213
rect 126532 3176 126560 3284
rect 127802 3272 127808 3324
rect 127860 3312 127866 3324
rect 128262 3312 128268 3324
rect 127860 3284 128268 3312
rect 127860 3272 127866 3284
rect 128262 3272 128268 3284
rect 128320 3272 128326 3324
rect 130120 3312 130148 3352
rect 150342 3340 150348 3392
rect 150400 3380 150406 3392
rect 155972 3380 156000 3420
rect 482278 3408 482284 3420
rect 482336 3408 482342 3460
rect 482370 3408 482376 3460
rect 482428 3448 482434 3460
rect 496538 3448 496544 3460
rect 482428 3420 496544 3448
rect 482428 3408 482434 3420
rect 496538 3408 496544 3420
rect 496596 3408 496602 3460
rect 497458 3408 497464 3460
rect 497516 3448 497522 3460
rect 509602 3448 509608 3460
rect 497516 3420 509608 3448
rect 497516 3408 497522 3420
rect 509602 3408 509608 3420
rect 509660 3408 509666 3460
rect 514570 3408 514576 3460
rect 514628 3448 514634 3460
rect 577406 3448 577412 3460
rect 514628 3420 577412 3448
rect 514628 3408 514634 3420
rect 577406 3408 577412 3420
rect 577464 3408 577470 3460
rect 150400 3352 156000 3380
rect 150400 3340 150406 3352
rect 156322 3340 156328 3392
rect 156380 3380 156386 3392
rect 157242 3380 157248 3392
rect 156380 3352 157248 3380
rect 156380 3340 156386 3352
rect 157242 3340 157248 3352
rect 157300 3340 157306 3392
rect 157518 3340 157524 3392
rect 157576 3380 157582 3392
rect 158622 3380 158628 3392
rect 157576 3352 158628 3380
rect 157576 3340 157582 3352
rect 158622 3340 158628 3352
rect 158680 3340 158686 3392
rect 158714 3340 158720 3392
rect 158772 3380 158778 3392
rect 160002 3380 160008 3392
rect 158772 3352 160008 3380
rect 158772 3340 158778 3352
rect 160002 3340 160008 3352
rect 160060 3340 160066 3392
rect 175366 3340 175372 3392
rect 175424 3380 175430 3392
rect 176562 3380 176568 3392
rect 175424 3352 176568 3380
rect 175424 3340 175430 3352
rect 176562 3340 176568 3352
rect 176620 3340 176626 3392
rect 181346 3340 181352 3392
rect 181404 3380 181410 3392
rect 182082 3380 182088 3392
rect 181404 3352 182088 3380
rect 181404 3340 181410 3352
rect 182082 3340 182088 3352
rect 182140 3340 182146 3392
rect 183554 3340 183560 3392
rect 183612 3380 183618 3392
rect 184842 3380 184848 3392
rect 183612 3352 184848 3380
rect 183612 3340 183618 3352
rect 184842 3340 184848 3352
rect 184900 3340 184906 3392
rect 231302 3340 231308 3392
rect 231360 3380 231366 3392
rect 231762 3380 231768 3392
rect 231360 3352 231768 3380
rect 231360 3340 231366 3352
rect 231762 3340 231768 3352
rect 231820 3340 231826 3392
rect 252554 3340 252560 3392
rect 252612 3380 252618 3392
rect 253842 3380 253848 3392
rect 252612 3352 253848 3380
rect 252612 3340 252618 3352
rect 253842 3340 253848 3352
rect 253900 3340 253906 3392
rect 261018 3340 261024 3392
rect 261076 3380 261082 3392
rect 262122 3380 262128 3392
rect 261076 3352 262128 3380
rect 261076 3340 261082 3352
rect 262122 3340 262128 3352
rect 262180 3340 262186 3392
rect 262214 3340 262220 3392
rect 262272 3380 262278 3392
rect 263502 3380 263508 3392
rect 262272 3352 263508 3380
rect 262272 3340 262278 3352
rect 263502 3340 263508 3352
rect 263560 3340 263566 3392
rect 263597 3383 263655 3389
rect 263597 3349 263609 3383
rect 263643 3380 263655 3383
rect 285674 3380 285680 3392
rect 263643 3352 285680 3380
rect 263643 3349 263655 3352
rect 263597 3343 263655 3349
rect 285674 3340 285680 3352
rect 285732 3340 285738 3392
rect 287054 3340 287060 3392
rect 287112 3380 287118 3392
rect 288342 3380 288348 3392
rect 287112 3352 288348 3380
rect 287112 3340 287118 3352
rect 288342 3340 288348 3352
rect 288400 3340 288406 3392
rect 296714 3340 296720 3392
rect 296772 3380 296778 3392
rect 297910 3380 297916 3392
rect 296772 3352 297916 3380
rect 296772 3340 296778 3352
rect 297910 3340 297916 3352
rect 297968 3340 297974 3392
rect 313274 3340 313280 3392
rect 313332 3380 313338 3392
rect 314562 3380 314568 3392
rect 313332 3352 314568 3380
rect 313332 3340 313338 3352
rect 314562 3340 314568 3352
rect 314620 3340 314626 3392
rect 321554 3340 321560 3392
rect 321612 3380 321618 3392
rect 322842 3380 322848 3392
rect 321612 3352 322848 3380
rect 321612 3340 321618 3352
rect 322842 3340 322848 3352
rect 322900 3340 322906 3392
rect 347774 3340 347780 3392
rect 347832 3380 347838 3392
rect 349062 3380 349068 3392
rect 347832 3352 349068 3380
rect 347832 3340 347838 3352
rect 349062 3340 349068 3352
rect 349120 3340 349126 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 366910 3380 366916 3392
rect 365772 3352 366916 3380
rect 365772 3340 365778 3352
rect 366910 3340 366916 3352
rect 366968 3340 366974 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375190 3380 375196 3392
rect 374052 3352 375196 3380
rect 374052 3340 374058 3352
rect 375190 3340 375196 3352
rect 375248 3340 375254 3392
rect 425057 3383 425115 3389
rect 425057 3349 425069 3383
rect 425103 3380 425115 3383
rect 428734 3380 428740 3392
rect 425103 3352 428740 3380
rect 425103 3349 425115 3352
rect 425057 3343 425115 3349
rect 428734 3340 428740 3352
rect 428792 3340 428798 3392
rect 442994 3340 443000 3392
rect 443052 3380 443058 3392
rect 444190 3380 444196 3392
rect 443052 3352 444196 3380
rect 443052 3340 443058 3352
rect 444190 3340 444196 3352
rect 444248 3340 444254 3392
rect 467926 3340 467932 3392
rect 467984 3380 467990 3392
rect 469122 3380 469128 3392
rect 467984 3352 469128 3380
rect 467984 3340 467990 3352
rect 469122 3340 469128 3352
rect 469180 3340 469186 3392
rect 150434 3312 150440 3324
rect 130120 3284 150440 3312
rect 150434 3272 150440 3284
rect 150492 3272 150498 3324
rect 240778 3272 240784 3324
rect 240836 3312 240842 3324
rect 241422 3312 241428 3324
rect 240836 3284 241428 3312
rect 240836 3272 240842 3284
rect 241422 3272 241428 3284
rect 241480 3272 241486 3324
rect 259822 3272 259828 3324
rect 259880 3312 259886 3324
rect 285858 3312 285864 3324
rect 259880 3284 285864 3312
rect 259880 3272 259886 3284
rect 285858 3272 285864 3284
rect 285916 3272 285922 3324
rect 128357 3247 128415 3253
rect 128357 3213 128369 3247
rect 128403 3244 128415 3247
rect 142062 3244 142068 3256
rect 128403 3216 142068 3244
rect 128403 3213 128415 3216
rect 128357 3207 128415 3213
rect 142062 3204 142068 3216
rect 142120 3204 142126 3256
rect 268102 3204 268108 3256
rect 268160 3244 268166 3256
rect 269022 3244 269028 3256
rect 268160 3216 269028 3244
rect 268160 3204 268166 3216
rect 269022 3204 269028 3216
rect 269080 3204 269086 3256
rect 276474 3204 276480 3256
rect 276532 3244 276538 3256
rect 281534 3244 281540 3256
rect 276532 3216 281540 3244
rect 276532 3204 276538 3216
rect 281534 3204 281540 3216
rect 281592 3204 281598 3256
rect 130194 3176 130200 3188
rect 126532 3148 130200 3176
rect 130194 3136 130200 3148
rect 130252 3136 130258 3188
rect 258626 3136 258632 3188
rect 258684 3176 258690 3188
rect 263597 3179 263655 3185
rect 263597 3176 263609 3179
rect 258684 3148 263609 3176
rect 258684 3136 258690 3148
rect 263597 3145 263609 3148
rect 263643 3145 263655 3179
rect 263597 3139 263655 3145
rect 94501 3111 94559 3117
rect 94501 3077 94513 3111
rect 94547 3108 94559 3111
rect 104161 3111 104219 3117
rect 104161 3108 104173 3111
rect 94547 3080 104173 3108
rect 94547 3077 94559 3080
rect 94501 3071 94559 3077
rect 104161 3077 104173 3080
rect 104207 3077 104219 3111
rect 104161 3071 104219 3077
rect 113652 3080 122880 3108
rect 99190 3000 99196 3052
rect 99248 3040 99254 3052
rect 113652 3040 113680 3080
rect 99248 3012 113680 3040
rect 113729 3043 113787 3049
rect 99248 3000 99254 3012
rect 113729 3009 113741 3043
rect 113775 3040 113787 3043
rect 122742 3040 122748 3052
rect 113775 3012 122748 3040
rect 113775 3009 113787 3012
rect 113729 3003 113787 3009
rect 122742 3000 122748 3012
rect 122800 3000 122806 3052
rect 122852 3040 122880 3080
rect 132586 3040 132592 3052
rect 122852 3012 132592 3040
rect 132586 3000 132592 3012
rect 132644 3000 132650 3052
rect 207474 3000 207480 3052
rect 207532 3040 207538 3052
rect 208302 3040 208308 3052
rect 207532 3012 208308 3040
rect 207532 3000 207538 3012
rect 208302 3000 208308 3012
rect 208360 3000 208366 3052
rect 165890 2932 165896 2984
rect 165948 2972 165954 2984
rect 166902 2972 166908 2984
rect 165948 2944 166908 2972
rect 165948 2932 165954 2944
rect 166902 2932 166908 2944
rect 166960 2932 166966 2984
rect 106277 2907 106335 2913
rect 106277 2873 106289 2907
rect 106323 2904 106335 2907
rect 113729 2907 113787 2913
rect 113729 2904 113741 2907
rect 106323 2876 113741 2904
rect 106323 2873 106335 2876
rect 106277 2867 106335 2873
rect 113729 2873 113741 2876
rect 113775 2873 113787 2907
rect 113729 2867 113787 2873
rect 193214 2864 193220 2916
rect 193272 2904 193278 2916
rect 194410 2904 194416 2916
rect 193272 2876 194416 2904
rect 193272 2864 193278 2876
rect 194410 2864 194416 2876
rect 194468 2864 194474 2916
rect 152737 2839 152795 2845
rect 152737 2805 152749 2839
rect 152783 2836 152795 2839
rect 153102 2836 153108 2848
rect 152783 2808 153108 2836
rect 152783 2805 152795 2808
rect 152737 2799 152795 2805
rect 153102 2796 153108 2808
rect 153160 2796 153166 2848
rect 194502 2836 194508 2848
rect 193232 2808 194508 2836
rect 193232 2780 193260 2808
rect 194502 2796 194508 2808
rect 194560 2796 194566 2848
rect 280062 2796 280068 2848
rect 280120 2836 280126 2848
rect 490558 2836 490564 2848
rect 280120 2808 490564 2836
rect 280120 2796 280126 2808
rect 490558 2796 490564 2808
rect 490616 2796 490622 2848
rect 193214 2728 193220 2780
rect 193272 2728 193278 2780
rect 152734 592 152740 604
rect 152695 564 152740 592
rect 152734 552 152740 564
rect 152792 552 152798 604
rect 186314 552 186320 604
rect 186372 592 186378 604
rect 187234 592 187240 604
rect 186372 564 187240 592
rect 186372 552 186378 564
rect 187234 552 187240 564
rect 187292 552 187298 604
rect 187694 552 187700 604
rect 187752 592 187758 604
rect 188430 592 188436 604
rect 187752 564 188436 592
rect 187752 552 187758 564
rect 188430 552 188436 564
rect 188488 552 188494 604
rect 236086 552 236092 604
rect 236144 592 236150 604
rect 237190 592 237196 604
rect 236144 564 237196 592
rect 236144 552 236150 564
rect 237190 552 237196 564
rect 237248 552 237254 604
rect 237558 552 237564 604
rect 237616 592 237622 604
rect 238386 592 238392 604
rect 237616 564 238392 592
rect 237616 552 237622 564
rect 238386 552 238392 564
rect 238444 552 238450 604
rect 280154 552 280160 604
rect 280212 592 280218 604
rect 281258 592 281264 604
rect 280212 564 281264 592
rect 280212 552 280218 564
rect 281258 552 281264 564
rect 281316 552 281322 604
rect 316034 552 316040 604
rect 316092 592 316098 604
rect 316954 592 316960 604
rect 316092 564 316960 592
rect 316092 552 316098 564
rect 316954 552 316960 564
rect 317012 552 317018 604
rect 318794 552 318800 604
rect 318852 592 318858 604
rect 319254 592 319260 604
rect 318852 564 319260 592
rect 318852 552 318858 564
rect 319254 552 319260 564
rect 319312 552 319318 604
rect 322934 552 322940 604
rect 322992 592 322998 604
rect 324038 592 324044 604
rect 322992 564 324044 592
rect 322992 552 322998 564
rect 324038 552 324044 564
rect 324096 552 324102 604
rect 324314 552 324320 604
rect 324372 592 324378 604
rect 325234 592 325240 604
rect 324372 564 325240 592
rect 324372 552 324378 564
rect 325234 552 325240 564
rect 325292 552 325298 604
rect 393314 552 393320 604
rect 393372 592 393378 604
rect 394234 592 394240 604
rect 393372 564 394240 592
rect 393372 552 393378 564
rect 394234 552 394240 564
rect 394292 552 394298 604
rect 396074 552 396080 604
rect 396132 592 396138 604
rect 396626 592 396632 604
rect 396132 564 396632 592
rect 396132 552 396138 564
rect 396626 552 396632 564
rect 396684 552 396690 604
rect 401594 552 401600 604
rect 401652 592 401658 604
rect 402514 592 402520 604
rect 401652 564 402520 592
rect 401652 552 401658 564
rect 402514 552 402520 564
rect 402572 552 402578 604
rect 412634 552 412640 604
rect 412692 592 412698 604
rect 413278 592 413284 604
rect 412692 564 413284 592
rect 412692 552 412698 564
rect 413278 552 413284 564
rect 413336 552 413342 604
rect 415394 552 415400 604
rect 415452 592 415458 604
rect 415670 592 415676 604
rect 415452 564 415676 592
rect 415452 552 415458 564
rect 415670 552 415676 564
rect 415728 552 415734 604
rect 418154 552 418160 604
rect 418212 592 418218 604
rect 419166 592 419172 604
rect 418212 564 419172 592
rect 418212 552 418218 564
rect 419166 552 419172 564
rect 419224 552 419230 604
rect 419534 552 419540 604
rect 419592 592 419598 604
rect 420362 592 420368 604
rect 419592 564 420368 592
rect 419592 552 419598 564
rect 420362 552 420368 564
rect 420420 552 420426 604
rect 547874 552 547880 604
rect 547932 592 547938 604
rect 548886 592 548892 604
rect 547932 564 548892 592
rect 547932 552 547938 564
rect 548886 552 548892 564
rect 548944 552 548950 604
rect 549254 552 549260 604
rect 549312 592 549318 604
rect 550082 592 550088 604
rect 549312 564 550088 592
rect 549312 552 549318 564
rect 550082 552 550088 564
rect 550140 552 550146 604
rect 556154 552 556160 604
rect 556212 592 556218 604
rect 557166 592 557172 604
rect 556212 564 557172 592
rect 556212 552 556218 564
rect 557166 552 557172 564
rect 557224 552 557230 604
rect 581086 552 581092 604
rect 581144 592 581150 604
rect 582190 592 582196 604
rect 581144 564 582196 592
rect 581144 552 581150 564
rect 582190 552 582196 564
rect 582248 552 582254 604
<< via1 >>
rect 111708 700680 111760 700732
rect 154120 700680 154172 700732
rect 105452 700612 105504 700664
rect 169760 700612 169812 700664
rect 235172 700612 235224 700664
rect 235908 700612 235960 700664
rect 137836 700544 137888 700596
rect 283012 700544 283064 700596
rect 72976 700476 73028 700528
rect 269120 700476 269172 700528
rect 287704 700476 287756 700528
rect 332508 700476 332560 700528
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 143448 700408 143500 700460
rect 348792 700408 348844 700460
rect 24308 700340 24360 700392
rect 253940 700340 253992 700392
rect 290464 700340 290516 700392
rect 413652 700340 413704 700392
rect 104808 700272 104860 700324
rect 397460 700272 397512 700324
rect 399484 700272 399536 700324
rect 478512 700272 478564 700324
rect 533344 700272 533396 700324
rect 559656 700272 559708 700324
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 542728 698232 542780 698284
rect 543556 698232 543608 698284
rect 319444 696940 319496 696992
rect 580172 696940 580224 696992
rect 8208 695444 8260 695496
rect 282920 692792 282972 692844
rect 283840 692792 283892 692844
rect 542728 688644 542780 688696
rect 299664 688576 299716 688628
rect 300124 688576 300176 688628
rect 429384 688576 429436 688628
rect 429844 688576 429896 688628
rect 542544 688576 542596 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 295984 685856 296036 685908
rect 580172 685856 580224 685908
rect 299572 684428 299624 684480
rect 429292 684428 429344 684480
rect 542452 684428 542504 684480
rect 3332 681708 3384 681760
rect 4804 681708 4856 681760
rect 8116 678988 8168 679040
rect 8024 678920 8076 678972
rect 364340 676175 364392 676184
rect 364340 676141 364349 676175
rect 364349 676141 364383 676175
rect 364383 676141 364392 676175
rect 364340 676132 364392 676141
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 60648 673480 60700 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 51724 667904 51776 667956
rect 299940 666544 299992 666596
rect 364432 666544 364484 666596
rect 429660 666544 429712 666596
rect 494152 666544 494204 666596
rect 542820 666544 542872 666596
rect 8024 654100 8076 654152
rect 8208 654100 8260 654152
rect 364340 654100 364392 654152
rect 364524 654100 364576 654152
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 313924 650020 313976 650072
rect 580172 650020 580224 650072
rect 299664 647232 299716 647284
rect 299756 647232 299808 647284
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 542544 647232 542596 647284
rect 542636 647232 542688 647284
rect 299664 640364 299716 640416
rect 299756 640364 299808 640416
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 542544 640364 542596 640416
rect 542636 640364 542688 640416
rect 293224 638936 293276 638988
rect 580172 638936 580224 638988
rect 8024 634788 8076 634840
rect 8208 634788 8260 634840
rect 364340 634788 364392 634840
rect 364524 634788 364576 634840
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 299572 630640 299624 630692
rect 299756 630640 299808 630692
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 542452 630640 542504 630692
rect 542636 630640 542688 630692
rect 284944 626560 284996 626612
rect 580172 626560 580224 626612
rect 4068 623772 4120 623824
rect 6184 623772 6236 623824
rect 8024 615476 8076 615528
rect 8208 615476 8260 615528
rect 364340 615476 364392 615528
rect 364524 615476 364576 615528
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 299572 611328 299624 611380
rect 299756 611328 299808 611380
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 542452 611328 542504 611380
rect 542636 611328 542688 611380
rect 3424 609968 3476 610020
rect 14556 609968 14608 610020
rect 299664 608583 299716 608592
rect 299664 608549 299673 608583
rect 299673 608549 299707 608583
rect 299707 608549 299716 608583
rect 299664 608540 299716 608549
rect 429384 608583 429436 608592
rect 429384 608549 429393 608583
rect 429393 608549 429427 608583
rect 429427 608549 429436 608583
rect 429384 608540 429436 608549
rect 542544 608583 542596 608592
rect 542544 608549 542553 608583
rect 542553 608549 542587 608583
rect 542587 608549 542596 608583
rect 542544 608540 542596 608549
rect 223488 603100 223540 603152
rect 580172 603100 580224 603152
rect 299848 601672 299900 601724
rect 429568 601672 429620 601724
rect 542728 601672 542780 601724
rect 299848 598927 299900 598936
rect 299848 598893 299857 598927
rect 299857 598893 299891 598927
rect 299891 598893 299900 598927
rect 299848 598884 299900 598893
rect 429568 598927 429620 598936
rect 429568 598893 429577 598927
rect 429577 598893 429611 598927
rect 429611 598893 429620 598927
rect 429568 598884 429620 598893
rect 542728 598927 542780 598936
rect 542728 598893 542737 598927
rect 542737 598893 542771 598927
rect 542771 598893 542780 598927
rect 542728 598884 542780 598893
rect 8024 596164 8076 596216
rect 8208 596164 8260 596216
rect 364340 596164 364392 596216
rect 364524 596164 364576 596216
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3240 594804 3292 594856
rect 190460 594804 190512 594856
rect 73068 592016 73120 592068
rect 580172 592016 580224 592068
rect 299940 589296 299992 589348
rect 429660 589296 429712 589348
rect 542820 589296 542872 589348
rect 8024 589271 8076 589280
rect 8024 589237 8033 589271
rect 8033 589237 8067 589271
rect 8067 589237 8076 589271
rect 8024 589228 8076 589237
rect 364156 589228 364208 589280
rect 364432 589228 364484 589280
rect 493876 589228 493928 589280
rect 494152 589228 494204 589280
rect 299940 582428 299992 582480
rect 429660 582428 429712 582480
rect 542820 582428 542872 582480
rect 299848 582292 299900 582344
rect 429568 582292 429620 582344
rect 542728 582292 542780 582344
rect 8024 579751 8076 579760
rect 8024 579717 8033 579751
rect 8033 579717 8067 579751
rect 8067 579717 8076 579751
rect 8024 579708 8076 579717
rect 329104 579640 329156 579692
rect 580172 579640 580224 579692
rect 7932 579572 7984 579624
rect 8116 579572 8168 579624
rect 4068 567196 4120 567248
rect 255320 567196 255372 567248
rect 429292 563116 429344 563168
rect 542452 563116 542504 563168
rect 429292 562980 429344 563032
rect 542452 562980 542504 563032
rect 7932 562912 7984 562964
rect 8116 562912 8168 562964
rect 429292 560235 429344 560244
rect 429292 560201 429301 560235
rect 429301 560201 429335 560235
rect 429335 560201 429344 560235
rect 429292 560192 429344 560201
rect 542452 560235 542504 560244
rect 542452 560201 542461 560235
rect 542461 560201 542495 560235
rect 542495 560201 542504 560235
rect 542452 560192 542504 560201
rect 521660 556384 521712 556436
rect 529296 556384 529348 556436
rect 415400 556316 415452 556368
rect 424876 556316 424928 556368
rect 364524 553435 364576 553444
rect 364524 553401 364533 553435
rect 364533 553401 364567 553435
rect 364567 553401 364576 553435
rect 364524 553392 364576 553401
rect 494244 553435 494296 553444
rect 494244 553401 494253 553435
rect 494253 553401 494287 553435
rect 494287 553401 494296 553435
rect 494244 553392 494296 553401
rect 4068 552032 4120 552084
rect 15844 552032 15896 552084
rect 299480 550604 299532 550656
rect 299664 550604 299716 550656
rect 364524 550647 364576 550656
rect 364524 550613 364533 550647
rect 364533 550613 364567 550647
rect 364567 550613 364576 550647
rect 364524 550604 364576 550613
rect 429476 550604 429528 550656
rect 494244 550647 494296 550656
rect 494244 550613 494253 550647
rect 494253 550613 494287 550647
rect 494287 550613 494296 550647
rect 494244 550604 494296 550613
rect 542636 550604 542688 550656
rect 8024 550579 8076 550588
rect 8024 550545 8033 550579
rect 8033 550545 8067 550579
rect 8067 550545 8076 550579
rect 8024 550536 8076 550545
rect 281448 545096 281500 545148
rect 580172 545096 580224 545148
rect 364524 543804 364576 543856
rect 494244 543804 494296 543856
rect 364616 543736 364668 543788
rect 494336 543736 494388 543788
rect 299296 543668 299348 543720
rect 299480 543668 299532 543720
rect 429292 543600 429344 543652
rect 429476 543600 429528 543652
rect 542452 543600 542504 543652
rect 542636 543600 542688 543652
rect 8208 540948 8260 541000
rect 3976 538432 4028 538484
rect 10324 538432 10376 538484
rect 429292 534012 429344 534064
rect 429476 534012 429528 534064
rect 542452 534012 542504 534064
rect 542636 534012 542688 534064
rect 249708 532720 249760 532772
rect 580172 532720 580224 532772
rect 299572 531292 299624 531344
rect 299756 531292 299808 531344
rect 364432 531292 364484 531344
rect 364708 531292 364760 531344
rect 494152 531292 494204 531344
rect 494428 531292 494480 531344
rect 299756 524424 299808 524476
rect 364708 524492 364760 524544
rect 429476 524424 429528 524476
rect 299848 524356 299900 524408
rect 364616 524356 364668 524408
rect 494428 524492 494480 524544
rect 542636 524424 542688 524476
rect 429568 524356 429620 524408
rect 494336 524356 494388 524408
rect 542728 524356 542780 524408
rect 8208 521636 8260 521688
rect 8392 521636 8444 521688
rect 299664 511980 299716 512032
rect 299940 511980 299992 512032
rect 364432 511980 364484 512032
rect 364708 511980 364760 512032
rect 429384 511980 429436 512032
rect 429660 511980 429712 512032
rect 494152 511980 494204 512032
rect 494428 511980 494480 512032
rect 542544 511980 542596 512032
rect 542820 511980 542872 512032
rect 3884 509260 3936 509312
rect 242900 509260 242952 509312
rect 285036 509260 285088 509312
rect 580172 509260 580224 509312
rect 8208 502324 8260 502376
rect 8392 502324 8444 502376
rect 299756 502324 299808 502376
rect 299940 502324 299992 502376
rect 364524 502324 364576 502376
rect 364708 502324 364760 502376
rect 429476 502324 429528 502376
rect 429660 502324 429712 502376
rect 494244 502324 494296 502376
rect 494428 502324 494480 502376
rect 542636 502324 542688 502376
rect 542820 502324 542872 502376
rect 294604 498176 294656 498228
rect 580172 498176 580224 498228
rect 4068 495456 4120 495508
rect 205640 495456 205692 495508
rect 7932 492600 7984 492652
rect 8116 492600 8168 492652
rect 299664 492643 299716 492652
rect 299664 492609 299673 492643
rect 299673 492609 299707 492643
rect 299707 492609 299716 492643
rect 299664 492600 299716 492609
rect 429384 492643 429436 492652
rect 429384 492609 429393 492643
rect 429393 492609 429427 492643
rect 429427 492609 429436 492643
rect 429384 492600 429436 492609
rect 542544 492643 542596 492652
rect 542544 492609 542553 492643
rect 542553 492609 542587 492643
rect 542587 492609 542596 492643
rect 542544 492600 542596 492609
rect 291844 485800 291896 485852
rect 580172 485800 580224 485852
rect 299664 485775 299716 485784
rect 299664 485741 299673 485775
rect 299673 485741 299707 485775
rect 299707 485741 299716 485775
rect 299664 485732 299716 485741
rect 429384 485775 429436 485784
rect 429384 485741 429393 485775
rect 429393 485741 429427 485775
rect 429427 485741 429436 485775
rect 429384 485732 429436 485741
rect 542544 485775 542596 485784
rect 542544 485741 542553 485775
rect 542553 485741 542587 485775
rect 542587 485741 542596 485775
rect 542544 485732 542596 485741
rect 3332 480564 3384 480616
rect 11704 480564 11756 480616
rect 364340 480224 364392 480276
rect 364524 480224 364576 480276
rect 494060 480224 494112 480276
rect 494244 480224 494296 480276
rect 299572 476076 299624 476128
rect 299756 476076 299808 476128
rect 429292 476076 429344 476128
rect 429476 476076 429528 476128
rect 542452 476076 542504 476128
rect 542636 476076 542688 476128
rect 8024 473288 8076 473340
rect 8116 473288 8168 473340
rect 299664 473331 299716 473340
rect 299664 473297 299673 473331
rect 299673 473297 299707 473331
rect 299707 473297 299716 473331
rect 299664 473288 299716 473297
rect 429384 473331 429436 473340
rect 429384 473297 429393 473331
rect 429393 473297 429427 473331
rect 429427 473297 429436 473331
rect 429384 473288 429436 473297
rect 542544 473331 542596 473340
rect 542544 473297 542553 473331
rect 542553 473297 542587 473331
rect 542587 473297 542596 473331
rect 542544 473288 542596 473297
rect 299664 466395 299716 466404
rect 299664 466361 299673 466395
rect 299673 466361 299707 466395
rect 299707 466361 299716 466395
rect 299664 466352 299716 466361
rect 429384 466395 429436 466404
rect 429384 466361 429393 466395
rect 429393 466361 429427 466395
rect 429427 466361 429436 466395
rect 429384 466352 429436 466361
rect 542544 466395 542596 466404
rect 542544 466361 542553 466395
rect 542553 466361 542587 466395
rect 542587 466361 542596 466395
rect 542544 466352 542596 466361
rect 160008 462340 160060 462392
rect 580172 462340 580224 462392
rect 235908 461592 235960 461644
rect 281540 461592 281592 461644
rect 364340 460912 364392 460964
rect 364524 460912 364576 460964
rect 494060 460912 494112 460964
rect 494244 460912 494296 460964
rect 299388 460844 299440 460896
rect 299756 460844 299808 460896
rect 100668 451256 100720 451308
rect 580172 451256 580224 451308
rect 299480 449871 299532 449880
rect 299480 449837 299489 449871
rect 299489 449837 299523 449871
rect 299523 449837 299532 449871
rect 299480 449828 299532 449837
rect 8024 447108 8076 447160
rect 429200 447108 429252 447160
rect 542360 447108 542412 447160
rect 8116 447040 8168 447092
rect 429292 447040 429344 447092
rect 542452 447040 542504 447092
rect 7840 444320 7892 444372
rect 8116 444320 8168 444372
rect 429016 444320 429068 444372
rect 429292 444320 429344 444372
rect 542176 444320 542228 444372
rect 542452 444320 542504 444372
rect 364340 441600 364392 441652
rect 364524 441600 364576 441652
rect 494060 441600 494112 441652
rect 494244 441600 494296 441652
rect 299572 440240 299624 440292
rect 62488 438880 62540 438932
rect 580172 438880 580224 438932
rect 3792 437452 3844 437504
rect 14464 437452 14516 437504
rect 299572 436772 299624 436824
rect 8024 427864 8076 427916
rect 429200 427796 429252 427848
rect 542360 427796 542412 427848
rect 8024 427728 8076 427780
rect 429292 427728 429344 427780
rect 542452 427728 542504 427780
rect 429016 425008 429068 425060
rect 429292 425008 429344 425060
rect 542176 425008 542228 425060
rect 542452 425008 542504 425060
rect 4068 423648 4120 423700
rect 13084 423648 13136 423700
rect 299572 423648 299624 423700
rect 364340 422288 364392 422340
rect 364524 422288 364576 422340
rect 494060 422288 494112 422340
rect 494244 422288 494296 422340
rect 299572 422220 299624 422272
rect 299756 422220 299808 422272
rect 8024 418140 8076 418192
rect 8208 418140 8260 418192
rect 315304 415420 315356 415472
rect 580172 415420 580224 415472
rect 299480 412564 299532 412616
rect 299572 412564 299624 412616
rect 429200 408484 429252 408536
rect 542360 408484 542412 408536
rect 429292 408348 429344 408400
rect 542452 408348 542504 408400
rect 429292 405671 429344 405680
rect 429292 405637 429301 405671
rect 429301 405637 429335 405671
rect 429335 405637 429344 405671
rect 429292 405628 429344 405637
rect 542452 405671 542504 405680
rect 542452 405637 542461 405671
rect 542461 405637 542495 405671
rect 542495 405637 542504 405671
rect 542452 405628 542504 405637
rect 286324 404336 286376 404388
rect 580172 404336 580224 404388
rect 364340 402976 364392 403028
rect 364524 402976 364576 403028
rect 494060 402976 494112 403028
rect 494244 402976 494296 403028
rect 299204 401548 299256 401600
rect 299572 401548 299624 401600
rect 8024 398939 8076 398948
rect 8024 398905 8033 398939
rect 8033 398905 8067 398939
rect 8067 398905 8076 398939
rect 8024 398896 8076 398905
rect 429292 398803 429344 398812
rect 429292 398769 429301 398803
rect 429301 398769 429335 398803
rect 429335 398769 429344 398803
rect 429292 398760 429344 398769
rect 542452 398803 542504 398812
rect 542452 398769 542461 398803
rect 542461 398769 542495 398803
rect 542495 398769 542504 398803
rect 542452 398760 542504 398769
rect 4068 394680 4120 394732
rect 281632 394680 281684 394732
rect 286416 391960 286468 392012
rect 580172 391960 580224 392012
rect 299388 391892 299440 391944
rect 8024 390575 8076 390584
rect 8024 390541 8033 390575
rect 8033 390541 8067 390575
rect 8067 390541 8076 390575
rect 8024 390532 8076 390541
rect 429292 389172 429344 389224
rect 542452 389172 542504 389224
rect 299572 389079 299624 389088
rect 299572 389045 299581 389079
rect 299581 389045 299615 389079
rect 299615 389045 299624 389079
rect 299572 389036 299624 389045
rect 429292 389036 429344 389088
rect 542452 389036 542504 389088
rect 364340 383664 364392 383716
rect 364524 383664 364576 383716
rect 494060 383664 494112 383716
rect 494244 383664 494296 383716
rect 7840 380876 7892 380928
rect 8024 380876 8076 380928
rect 3976 379516 4028 379568
rect 24124 379516 24176 379568
rect 299572 379448 299624 379500
rect 299756 379448 299808 379500
rect 429292 379448 429344 379500
rect 429476 379448 429528 379500
rect 542452 379448 542504 379500
rect 542636 379448 542688 379500
rect 8024 369860 8076 369912
rect 7932 369792 7984 369844
rect 60556 368500 60608 368552
rect 580172 368500 580224 368552
rect 4068 365712 4120 365764
rect 183560 365712 183612 365764
rect 364524 360247 364576 360256
rect 364524 360213 364533 360247
rect 364533 360213 364567 360247
rect 364567 360213 364576 360247
rect 364524 360204 364576 360213
rect 494244 360247 494296 360256
rect 494244 360213 494253 360247
rect 494253 360213 494287 360247
rect 494287 360213 494296 360247
rect 494244 360204 494296 360213
rect 7932 360136 7984 360188
rect 8116 360136 8168 360188
rect 299848 357527 299900 357536
rect 299848 357493 299857 357527
rect 299857 357493 299891 357527
rect 299891 357493 299900 357527
rect 299848 357484 299900 357493
rect 364524 357527 364576 357536
rect 364524 357493 364533 357527
rect 364533 357493 364567 357527
rect 364567 357493 364576 357527
rect 364524 357484 364576 357493
rect 429568 357527 429620 357536
rect 429568 357493 429577 357527
rect 429577 357493 429611 357527
rect 429611 357493 429620 357527
rect 429568 357484 429620 357493
rect 494244 357527 494296 357536
rect 494244 357493 494253 357527
rect 494253 357493 494287 357527
rect 494287 357493 494296 357527
rect 494244 357484 494296 357493
rect 542728 357527 542780 357536
rect 542728 357493 542737 357527
rect 542737 357493 542771 357527
rect 542771 357493 542780 357527
rect 542728 357484 542780 357493
rect 304356 357416 304408 357468
rect 580172 357416 580224 357468
rect 8116 357348 8168 357400
rect 299756 356124 299808 356176
rect 299848 354671 299900 354680
rect 299848 354637 299857 354671
rect 299857 354637 299891 354671
rect 299891 354637 299900 354671
rect 299848 354628 299900 354637
rect 429568 353379 429620 353388
rect 429568 353345 429577 353379
rect 429577 353345 429611 353379
rect 429611 353345 429620 353379
rect 429568 353336 429620 353345
rect 542728 353379 542780 353388
rect 542728 353345 542737 353379
rect 542737 353345 542771 353379
rect 542771 353345 542780 353379
rect 542728 353336 542780 353345
rect 429660 353243 429712 353252
rect 429660 353209 429669 353243
rect 429669 353209 429703 353243
rect 429703 353209 429712 353243
rect 429660 353200 429712 353209
rect 542820 353243 542872 353252
rect 542820 353209 542829 353243
rect 542829 353209 542863 353243
rect 542863 353209 542872 353243
rect 542820 353200 542872 353209
rect 8024 347803 8076 347812
rect 8024 347769 8033 347803
rect 8033 347769 8067 347803
rect 8067 347769 8076 347803
rect 8024 347760 8076 347769
rect 364340 347735 364392 347744
rect 364340 347701 364349 347735
rect 364349 347701 364383 347735
rect 364383 347701 364392 347735
rect 364340 347692 364392 347701
rect 494060 347735 494112 347744
rect 494060 347701 494069 347735
rect 494069 347701 494103 347735
rect 494103 347701 494112 347735
rect 494060 347692 494112 347701
rect 285128 345040 285180 345092
rect 580172 345040 580224 345092
rect 8024 341003 8076 341012
rect 8024 340969 8033 341003
rect 8033 340969 8067 341003
rect 8067 340969 8076 341003
rect 8024 340960 8076 340969
rect 429660 340799 429712 340808
rect 429660 340765 429669 340799
rect 429669 340765 429703 340799
rect 429703 340765 429712 340799
rect 429660 340756 429712 340765
rect 542820 340799 542872 340808
rect 542820 340765 542829 340799
rect 542829 340765 542863 340799
rect 542863 340765 542872 340799
rect 542820 340756 542872 340765
rect 364432 338104 364484 338156
rect 494152 338104 494204 338156
rect 8024 336855 8076 336864
rect 8024 336821 8033 336855
rect 8033 336821 8067 336855
rect 8067 336821 8076 336855
rect 8024 336812 8076 336821
rect 4068 336744 4120 336796
rect 281908 336744 281960 336796
rect 299940 336744 299992 336796
rect 8024 336608 8076 336660
rect 7932 327131 7984 327140
rect 7932 327097 7941 327131
rect 7941 327097 7975 327131
rect 7975 327097 7984 327131
rect 7932 327088 7984 327097
rect 299756 327088 299808 327140
rect 299848 327088 299900 327140
rect 364340 325660 364392 325712
rect 364524 325660 364576 325712
rect 429476 325660 429528 325712
rect 429568 325660 429620 325712
rect 494060 325660 494112 325712
rect 494244 325660 494296 325712
rect 542636 325660 542688 325712
rect 542728 325660 542780 325712
rect 291936 321580 291988 321632
rect 580172 321580 580224 321632
rect 7932 321444 7984 321496
rect 8208 321444 8260 321496
rect 299664 318792 299716 318844
rect 299756 318792 299808 318844
rect 429384 318792 429436 318844
rect 429476 318792 429528 318844
rect 542544 318792 542596 318844
rect 542636 318792 542688 318844
rect 299664 311924 299716 311976
rect 299756 311924 299808 311976
rect 429384 311924 429436 311976
rect 429476 311924 429528 311976
rect 542544 311924 542596 311976
rect 542636 311924 542688 311976
rect 61200 310496 61252 310548
rect 579804 310496 579856 310548
rect 7932 309204 7984 309256
rect 8208 309204 8260 309256
rect 4068 307776 4120 307828
rect 22744 307776 22796 307828
rect 364340 306348 364392 306400
rect 364524 306348 364576 306400
rect 494060 306348 494112 306400
rect 494244 306348 494296 306400
rect 8024 302268 8076 302320
rect 299572 302200 299624 302252
rect 299756 302200 299808 302252
rect 429292 302200 429344 302252
rect 429476 302200 429528 302252
rect 542452 302200 542504 302252
rect 542636 302200 542688 302252
rect 8116 302064 8168 302116
rect 299664 299455 299716 299464
rect 299664 299421 299673 299455
rect 299673 299421 299707 299455
rect 299707 299421 299716 299455
rect 299664 299412 299716 299421
rect 216588 298120 216640 298172
rect 580172 298120 580224 298172
rect 3148 293972 3200 294024
rect 7564 293972 7616 294024
rect 299756 289824 299808 289876
rect 8208 289756 8260 289808
rect 429476 289799 429528 289808
rect 429476 289765 429485 289799
rect 429485 289765 429519 289799
rect 429519 289765 429528 289799
rect 429476 289756 429528 289765
rect 542636 289756 542688 289808
rect 364340 287036 364392 287088
rect 364524 287036 364576 287088
rect 494060 287036 494112 287088
rect 494244 287036 494296 287088
rect 286508 282140 286560 282192
rect 494060 282140 494112 282192
rect 8116 280211 8168 280220
rect 8116 280177 8125 280211
rect 8125 280177 8159 280211
rect 8159 280177 8168 280211
rect 8116 280168 8168 280177
rect 429568 280168 429620 280220
rect 542452 280211 542504 280220
rect 542452 280177 542461 280211
rect 542461 280177 542495 280211
rect 542495 280177 542504 280211
rect 542452 280168 542504 280177
rect 89628 277992 89680 278044
rect 283380 277992 283432 278044
rect 429384 274864 429436 274916
rect 429568 274864 429620 274916
rect 290556 274660 290608 274712
rect 580172 274660 580224 274712
rect 202788 273912 202840 273964
rect 283472 273912 283524 273964
rect 8116 273300 8168 273352
rect 8116 273096 8168 273148
rect 60464 272484 60516 272536
rect 462320 272484 462372 272536
rect 60924 271124 60976 271176
rect 527180 271124 527232 271176
rect 98644 270648 98696 270700
rect 443000 270648 443052 270700
rect 64052 270580 64104 270632
rect 458180 270580 458232 270632
rect 73804 270512 73856 270564
rect 476120 270512 476172 270564
rect 429384 270487 429436 270496
rect 429384 270453 429393 270487
rect 429393 270453 429427 270487
rect 429427 270453 429436 270487
rect 429384 270444 429436 270453
rect 97540 269968 97592 270020
rect 460940 269968 460992 270020
rect 120356 269900 120408 269952
rect 520280 269900 520332 269952
rect 189540 269832 189592 269884
rect 285956 269832 286008 269884
rect 22744 269764 22796 269816
rect 76748 269764 76800 269816
rect 187700 269764 187752 269816
rect 289820 269764 289872 269816
rect 164884 269696 164936 269748
rect 288532 269696 288584 269748
rect 156972 269628 157024 269680
rect 287152 269628 287204 269680
rect 152924 269560 152976 269612
rect 285680 269560 285732 269612
rect 181628 269492 181680 269544
rect 412640 269492 412692 269544
rect 174820 269424 174872 269476
rect 418160 269424 418212 269476
rect 139124 269356 139176 269408
rect 416872 269356 416924 269408
rect 163964 269288 164016 269340
rect 465080 269288 465132 269340
rect 112444 269220 112496 269272
rect 419540 269220 419592 269272
rect 262772 269152 262824 269204
rect 287244 269152 287296 269204
rect 260748 269084 260800 269136
rect 286048 269084 286100 269136
rect 163044 268608 163096 268660
rect 542452 268608 542504 268660
rect 220268 268540 220320 268592
rect 294696 268540 294748 268592
rect 211436 268472 211488 268524
rect 293316 268472 293368 268524
rect 172796 268404 172848 268456
rect 281816 268404 281868 268456
rect 178684 268336 178736 268388
rect 288624 268336 288676 268388
rect 213276 268268 213328 268320
rect 408500 268268 408552 268320
rect 55864 268200 55916 268252
rect 214380 268200 214432 268252
rect 236092 268200 236144 268252
rect 436100 268200 436152 268252
rect 69020 268132 69072 268184
rect 283288 268132 283340 268184
rect 6276 268064 6328 268116
rect 273628 268064 273680 268116
rect 168748 267996 168800 268048
rect 518900 267996 518952 268048
rect 19984 267928 20036 267980
rect 229100 267928 229152 267980
rect 230204 267928 230256 267980
rect 579804 267928 579856 267980
rect 188620 267860 188672 267912
rect 539600 267860 539652 267912
rect 145012 267792 145064 267844
rect 521660 267792 521712 267844
rect 252836 267724 252888 267776
rect 284392 267724 284444 267776
rect 542360 267724 542412 267776
rect 542636 267724 542688 267776
rect 99564 267656 99616 267708
rect 100668 267656 100720 267708
rect 110420 267656 110472 267708
rect 111708 267656 111760 267708
rect 248972 267656 249024 267708
rect 249708 267656 249760 267708
rect 280620 267656 280672 267708
rect 281448 267656 281500 267708
rect 89628 267316 89680 267368
rect 270500 267316 270552 267368
rect 259828 267248 259880 267300
rect 281356 267248 281408 267300
rect 115388 267180 115440 267232
rect 257988 267180 258040 267232
rect 263692 267180 263744 267232
rect 287888 267180 287940 267232
rect 249892 267112 249944 267164
rect 282276 267112 282328 267164
rect 84660 267044 84712 267096
rect 305000 267044 305052 267096
rect 57704 266976 57756 267028
rect 116308 266976 116360 267028
rect 265716 266976 265768 267028
rect 281172 266976 281224 267028
rect 57796 266908 57848 266960
rect 128268 266908 128320 266960
rect 132868 266908 132920 266960
rect 180708 266908 180760 266960
rect 237012 266908 237064 266960
rect 281724 266908 281776 266960
rect 57888 266840 57940 266892
rect 137100 266840 137152 266892
rect 226156 266840 226208 266892
rect 287796 266840 287848 266892
rect 56324 266772 56376 266824
rect 154948 266772 155000 266824
rect 164148 266772 164200 266824
rect 197452 266772 197504 266824
rect 198556 266772 198608 266824
rect 282000 266772 282052 266824
rect 56232 266704 56284 266756
rect 179788 266704 179840 266756
rect 194508 266704 194560 266756
rect 282460 266704 282512 266756
rect 67916 266636 67968 266688
rect 126980 266636 127032 266688
rect 256884 266636 256936 266688
rect 283104 266636 283156 266688
rect 17224 266568 17276 266620
rect 117412 266568 117464 266620
rect 124220 266568 124272 266620
rect 282368 266568 282420 266620
rect 157892 266500 157944 266552
rect 270684 266500 270736 266552
rect 283564 266500 283616 266552
rect 55128 266432 55180 266484
rect 66996 266432 67048 266484
rect 71964 266432 72016 266484
rect 259460 266432 259512 266484
rect 267740 266432 267792 266484
rect 288716 266432 288768 266484
rect 53748 266364 53800 266416
rect 65892 266364 65944 266416
rect 122380 266364 122432 266416
rect 128360 266364 128412 266416
rect 158996 266364 159048 266416
rect 160008 266364 160060 266416
rect 163412 266364 163464 266416
rect 210332 266364 210384 266416
rect 226248 266364 226300 266416
rect 277676 266364 277728 266416
rect 280896 266364 280948 266416
rect 3884 266296 3936 266348
rect 69020 266296 69072 266348
rect 263600 266339 263652 266348
rect 263600 266305 263609 266339
rect 263609 266305 263643 266339
rect 263643 266305 263652 266339
rect 263600 266296 263652 266305
rect 271788 266271 271840 266280
rect 271788 266237 271797 266271
rect 271797 266237 271831 266271
rect 271831 266237 271840 266271
rect 271788 266228 271840 266237
rect 155868 265820 155920 265872
rect 482284 265820 482336 265872
rect 231124 265752 231176 265804
rect 284300 265752 284352 265804
rect 3516 265684 3568 265736
rect 164148 265684 164200 265736
rect 257988 265684 258040 265736
rect 374000 265684 374052 265736
rect 128360 265616 128412 265668
rect 351920 265616 351972 265668
rect 275652 265548 275704 265600
rect 345020 265548 345072 265600
rect 215300 265480 215352 265532
rect 286140 265480 286192 265532
rect 221188 265412 221240 265464
rect 298100 265412 298152 265464
rect 149980 265344 150032 265396
rect 284576 265344 284628 265396
rect 96620 265276 96672 265328
rect 327080 265276 327132 265328
rect 171876 265208 171928 265260
rect 437480 265208 437532 265260
rect 161940 265140 161992 265192
rect 435364 265140 435416 265192
rect 68836 265072 68888 265124
rect 347780 265072 347832 265124
rect 233056 265004 233108 265056
rect 547880 265004 547932 265056
rect 268936 264936 268988 264988
rect 287060 264936 287112 264988
rect 285772 264596 285824 264648
rect 252192 264571 252244 264580
rect 252192 264537 252201 264571
rect 252201 264537 252235 264571
rect 252235 264537 252244 264571
rect 252192 264528 252244 264537
rect 259184 264571 259236 264580
rect 259184 264537 259193 264571
rect 259193 264537 259227 264571
rect 259227 264537 259236 264571
rect 259184 264528 259236 264537
rect 284668 264528 284720 264580
rect 161112 264460 161164 264512
rect 284484 264460 284536 264512
rect 81440 264299 81492 264308
rect 81440 264265 81449 264299
rect 81449 264265 81483 264299
rect 81483 264265 81492 264299
rect 81440 264256 81492 264265
rect 85580 264299 85632 264308
rect 85580 264265 85589 264299
rect 85589 264265 85623 264299
rect 85623 264265 85632 264299
rect 85580 264256 85632 264265
rect 87420 264299 87472 264308
rect 87420 264265 87429 264299
rect 87429 264265 87463 264299
rect 87463 264265 87472 264299
rect 87420 264256 87472 264265
rect 132868 264392 132920 264444
rect 208400 264392 208452 264444
rect 108672 264299 108724 264308
rect 108672 264265 108681 264299
rect 108681 264265 108715 264299
rect 108715 264265 108724 264299
rect 108672 264256 108724 264265
rect 136456 264324 136508 264376
rect 132316 264256 132368 264308
rect 133512 264299 133564 264308
rect 133512 264265 133521 264299
rect 133521 264265 133555 264299
rect 133555 264265 133564 264299
rect 133512 264256 133564 264265
rect 134432 264299 134484 264308
rect 134432 264265 134441 264299
rect 134441 264265 134475 264299
rect 134475 264265 134484 264299
rect 134432 264256 134484 264265
rect 144368 264256 144420 264308
rect 226248 264324 226300 264376
rect 242256 264324 242308 264376
rect 300860 264324 300912 264376
rect 147680 264299 147732 264308
rect 147680 264265 147689 264299
rect 147689 264265 147723 264299
rect 147723 264265 147732 264299
rect 147680 264256 147732 264265
rect 173808 264299 173860 264308
rect 173808 264265 173817 264299
rect 173817 264265 173851 264299
rect 173851 264265 173860 264299
rect 173808 264256 173860 264265
rect 202696 264299 202748 264308
rect 202696 264265 202705 264299
rect 202705 264265 202739 264299
rect 202739 264265 202748 264299
rect 202696 264256 202748 264265
rect 218520 264256 218572 264308
rect 224408 264299 224460 264308
rect 224408 264265 224417 264299
rect 224417 264265 224451 264299
rect 224451 264265 224460 264299
rect 224408 264256 224460 264265
rect 278688 264299 278740 264308
rect 278688 264265 278697 264299
rect 278697 264265 278731 264299
rect 278731 264265 278740 264299
rect 278688 264256 278740 264265
rect 279792 264256 279844 264308
rect 280804 264256 280856 264308
rect 492680 264188 492732 264240
rect 296720 264120 296772 264172
rect 498200 264052 498252 264104
rect 369860 263984 369912 264036
rect 361580 263916 361632 263968
rect 375380 263848 375432 263900
rect 56508 263780 56560 263832
rect 451280 263780 451332 263832
rect 56416 263712 56468 263764
rect 390560 263712 390612 263764
rect 55036 263644 55088 263696
rect 368480 263644 368532 263696
rect 53656 263576 53708 263628
rect 527180 263576 527232 263628
rect 281356 263508 281408 263560
rect 288440 263508 288492 263560
rect 429384 263551 429436 263560
rect 429384 263517 429393 263551
rect 429393 263517 429427 263551
rect 429427 263517 429436 263551
rect 429384 263508 429436 263517
rect 282184 263440 282236 263492
rect 282460 263440 282512 263492
rect 280988 263168 281040 263220
rect 556160 263168 556212 263220
rect 499580 263100 499632 263152
rect 285864 263032 285916 263084
rect 281080 262964 281132 263016
rect 357440 262896 357492 262948
rect 445760 262828 445812 262880
rect 60280 262760 60332 262812
rect 286600 262760 286652 262812
rect 282368 261604 282420 261656
rect 296812 261604 296864 261656
rect 281172 261536 281224 261588
rect 451372 261536 451424 261588
rect 280988 261468 281040 261520
rect 459560 261468 459612 261520
rect 1308 261400 1360 261452
rect 283196 260856 283248 260908
rect 304264 260856 304316 260908
rect 6184 260788 6236 260840
rect 59360 260788 59412 260840
rect 299480 260788 299532 260840
rect 299664 260788 299716 260840
rect 429384 260788 429436 260840
rect 280896 260176 280948 260228
rect 455420 260176 455472 260228
rect 281264 260108 281316 260160
rect 485780 260108 485832 260160
rect 283104 258748 283156 258800
rect 306380 258748 306432 258800
rect 282000 258680 282052 258732
rect 367100 258680 367152 258732
rect 282276 257320 282328 257372
rect 467840 257320 467892 257372
rect 283564 255960 283616 256012
rect 402980 255960 403032 256012
rect 429568 253963 429620 253972
rect 429568 253929 429577 253963
rect 429577 253929 429611 253963
rect 429611 253929 429620 253963
rect 429568 253920 429620 253929
rect 280804 253172 280856 253224
rect 578240 253172 578292 253224
rect 286600 252492 286652 252544
rect 579804 252492 579856 252544
rect 4068 251200 4120 251252
rect 8944 251200 8996 251252
rect 284116 251200 284168 251252
rect 332600 251200 332652 251252
rect 284208 251132 284260 251184
rect 304356 251132 304408 251184
rect 284208 248412 284260 248464
rect 302240 248412 302292 248464
rect 284208 245624 284260 245676
rect 311900 245624 311952 245676
rect 284208 244264 284260 244316
rect 535460 244264 535512 244316
rect 542360 244196 542412 244248
rect 542636 244196 542688 244248
rect 287980 243516 288032 243568
rect 400220 243516 400272 243568
rect 283840 238688 283892 238740
rect 319444 238688 319496 238740
rect 282184 238008 282236 238060
rect 396080 238008 396132 238060
rect 4068 237328 4120 237380
rect 17224 237328 17276 237380
rect 429292 234676 429344 234728
rect 429292 234540 429344 234592
rect 284208 233248 284260 233300
rect 308404 233248 308456 233300
rect 7932 231820 7984 231872
rect 8024 231820 8076 231872
rect 299480 231820 299532 231872
rect 299756 231820 299808 231872
rect 542544 231820 542596 231872
rect 542728 231820 542780 231872
rect 429292 231795 429344 231804
rect 429292 231761 429301 231795
rect 429301 231761 429335 231795
rect 429335 231761 429344 231795
rect 429292 231752 429344 231761
rect 284116 228556 284168 228608
rect 286508 228556 286560 228608
rect 284208 226312 284260 226364
rect 467104 226312 467156 226364
rect 284208 224952 284260 225004
rect 497464 224952 497516 225004
rect 3608 223524 3660 223576
rect 59360 223524 59412 223576
rect 2964 223456 3016 223508
rect 19984 223456 20036 223508
rect 429476 222164 429528 222216
rect 542360 222164 542412 222216
rect 542636 222164 542688 222216
rect 8024 222139 8076 222148
rect 8024 222105 8033 222139
rect 8033 222105 8067 222139
rect 8067 222105 8076 222139
rect 8024 222096 8076 222105
rect 53564 220804 53616 220856
rect 59360 220804 59412 220856
rect 53472 216656 53524 216708
rect 59452 216656 59504 216708
rect 284208 216656 284260 216708
rect 385684 216656 385736 216708
rect 14556 216588 14608 216640
rect 59360 216588 59412 216640
rect 284208 215296 284260 215348
rect 514024 215296 514076 215348
rect 8116 215160 8168 215212
rect 429292 215160 429344 215212
rect 429476 215160 429528 215212
rect 54944 213936 54996 213988
rect 59360 213936 59412 213988
rect 299480 212576 299532 212628
rect 299756 212576 299808 212628
rect 56140 212508 56192 212560
rect 59360 212508 59412 212560
rect 284208 212508 284260 212560
rect 331220 212508 331272 212560
rect 284208 211148 284260 211200
rect 462320 211148 462372 211200
rect 280896 209788 280948 209840
rect 281172 209788 281224 209840
rect 280804 209763 280856 209772
rect 280804 209729 280813 209763
rect 280813 209729 280847 209763
rect 280847 209729 280856 209763
rect 280804 209720 280856 209729
rect 284116 207000 284168 207052
rect 478880 207000 478932 207052
rect 8116 205708 8168 205760
rect 53380 205640 53432 205692
rect 59360 205640 59412 205692
rect 7932 205572 7984 205624
rect 429292 205572 429344 205624
rect 429476 205572 429528 205624
rect 284208 204348 284260 204400
rect 305644 204348 305696 204400
rect 304356 204280 304408 204332
rect 579896 204280 579948 204332
rect 54852 202852 54904 202904
rect 59360 202852 59412 202904
rect 542544 202852 542596 202904
rect 542636 202852 542688 202904
rect 299664 202827 299716 202836
rect 299664 202793 299673 202827
rect 299673 202793 299707 202827
rect 299707 202793 299716 202827
rect 299664 202784 299716 202793
rect 429476 202827 429528 202836
rect 429476 202793 429485 202827
rect 429485 202793 429519 202827
rect 429519 202793 429528 202827
rect 429476 202784 429528 202793
rect 284208 201492 284260 201544
rect 337384 201492 337436 201544
rect 7932 201467 7984 201476
rect 7932 201433 7941 201467
rect 7941 201433 7975 201467
rect 7975 201433 7984 201467
rect 7932 201424 7984 201433
rect 280988 200132 281040 200184
rect 24124 200064 24176 200116
rect 59360 200064 59412 200116
rect 280988 200039 281040 200048
rect 280988 200005 280997 200039
rect 280997 200005 281031 200039
rect 281031 200005 281040 200039
rect 280988 199996 281040 200005
rect 284208 198704 284260 198756
rect 430580 198704 430632 198756
rect 542636 195984 542688 196036
rect 542728 195916 542780 195968
rect 27620 194488 27672 194540
rect 37188 194488 37240 194540
rect 299756 193264 299808 193316
rect 429568 193264 429620 193316
rect 53288 193196 53340 193248
rect 59360 193196 59412 193248
rect 284208 193196 284260 193248
rect 517520 193196 517572 193248
rect 7932 193171 7984 193180
rect 7932 193137 7941 193171
rect 7941 193137 7975 193171
rect 7975 193137 7984 193171
rect 7932 193128 7984 193137
rect 280988 190859 281040 190868
rect 280988 190825 280997 190859
rect 280997 190825 281031 190859
rect 281031 190825 281040 190859
rect 280988 190816 281040 190825
rect 3700 188980 3752 189032
rect 59360 188980 59412 189032
rect 284208 187688 284260 187740
rect 364984 187688 365036 187740
rect 8024 186328 8076 186380
rect 8116 186192 8168 186244
rect 542544 183540 542596 183592
rect 542820 183540 542872 183592
rect 429476 183515 429528 183524
rect 429476 183481 429485 183515
rect 429485 183481 429519 183515
rect 429519 183481 429528 183515
rect 429476 183472 429528 183481
rect 57612 182180 57664 182232
rect 59912 182180 59964 182232
rect 284208 182180 284260 182232
rect 292580 182180 292632 182232
rect 293316 182112 293368 182164
rect 580172 182112 580224 182164
rect 53196 180820 53248 180872
rect 59360 180820 59412 180872
rect 280988 179324 281040 179376
rect 281448 179324 281500 179376
rect 8116 176740 8168 176792
rect 8024 176536 8076 176588
rect 284208 176672 284260 176724
rect 502984 176672 503036 176724
rect 57520 175244 57572 175296
rect 59544 175244 59596 175296
rect 299480 173952 299532 174004
rect 299756 173952 299808 174004
rect 429568 173952 429620 174004
rect 284208 173884 284260 173936
rect 477500 173884 477552 173936
rect 542636 173884 542688 173936
rect 542820 173884 542872 173936
rect 280804 171912 280856 171964
rect 281172 171912 281224 171964
rect 284208 171096 284260 171148
rect 447140 171096 447192 171148
rect 285312 169736 285364 169788
rect 580172 169736 580224 169788
rect 542360 169056 542412 169108
rect 542636 169056 542688 169108
rect 15844 168308 15896 168360
rect 59360 168308 59412 168360
rect 281264 166880 281316 166932
rect 281448 166880 281500 166932
rect 3332 165520 3384 165572
rect 6276 165520 6328 165572
rect 13084 165520 13136 165572
rect 59360 165520 59412 165572
rect 283840 164228 283892 164280
rect 501604 164228 501656 164280
rect 8024 164160 8076 164212
rect 8116 164160 8168 164212
rect 299480 164160 299532 164212
rect 299664 164160 299716 164212
rect 429384 164203 429436 164212
rect 429384 164169 429393 164203
rect 429393 164169 429427 164203
rect 429427 164169 429436 164203
rect 429384 164160 429436 164169
rect 283840 162868 283892 162920
rect 371884 162868 371936 162920
rect 280804 162120 280856 162172
rect 281264 162120 281316 162172
rect 542360 161372 542412 161424
rect 542636 161372 542688 161424
rect 283380 160080 283432 160132
rect 316040 160080 316092 160132
rect 422944 157360 422996 157412
rect 579896 157360 579948 157412
rect 429384 157335 429436 157344
rect 429384 157301 429393 157335
rect 429393 157301 429427 157335
rect 429427 157301 429436 157335
rect 429384 157292 429436 157301
rect 284024 153212 284076 153264
rect 322296 153212 322348 153264
rect 280804 152600 280856 152652
rect 281172 152600 281224 152652
rect 280804 152396 280856 152448
rect 281264 152396 281316 152448
rect 542360 151784 542412 151836
rect 542636 151784 542688 151836
rect 6184 150424 6236 150476
rect 59360 150424 59412 150476
rect 283840 150356 283892 150408
rect 315304 150356 315356 150408
rect 429292 147636 429344 147688
rect 429476 147636 429528 147688
rect 8024 144848 8076 144900
rect 8116 144848 8168 144900
rect 283840 144848 283892 144900
rect 422944 144848 422996 144900
rect 429384 144891 429436 144900
rect 429384 144857 429393 144891
rect 429393 144857 429427 144891
rect 429427 144857 429436 144891
rect 429384 144848 429436 144857
rect 57428 142604 57480 142656
rect 59360 142604 59412 142656
rect 283840 142128 283892 142180
rect 372620 142128 372672 142180
rect 284208 142060 284260 142112
rect 313924 142060 313976 142112
rect 542360 142060 542412 142112
rect 542636 142060 542688 142112
rect 429384 137955 429436 137964
rect 429384 137921 429393 137955
rect 429393 137921 429427 137955
rect 429427 137921 429436 137955
rect 429384 137912 429436 137921
rect 283748 136620 283800 136672
rect 426440 136620 426492 136672
rect 3976 135260 4028 135312
rect 53104 135260 53156 135312
rect 284208 135260 284260 135312
rect 354680 135260 354732 135312
rect 280988 135192 281040 135244
rect 308496 133900 308548 133952
rect 580172 133900 580224 133952
rect 542360 132472 542412 132524
rect 542636 132472 542688 132524
rect 58532 131112 58584 131164
rect 59360 131112 59412 131164
rect 57244 129752 57296 129804
rect 59728 129752 59780 129804
rect 54760 128324 54812 128376
rect 59360 128324 59412 128376
rect 60648 128324 60700 128376
rect 62396 128324 62448 128376
rect 429292 128324 429344 128376
rect 429476 128324 429528 128376
rect 542360 128256 542412 128308
rect 542636 128256 542688 128308
rect 282184 127576 282236 127628
rect 283564 127576 283616 127628
rect 280896 125715 280948 125724
rect 280896 125681 280905 125715
rect 280905 125681 280939 125715
rect 280939 125681 280948 125715
rect 280896 125672 280948 125681
rect 8024 125536 8076 125588
rect 280896 125579 280948 125588
rect 280896 125545 280905 125579
rect 280905 125545 280939 125579
rect 280939 125545 280948 125579
rect 280896 125536 280948 125545
rect 429292 125579 429344 125588
rect 429292 125545 429301 125579
rect 429301 125545 429335 125579
rect 429335 125545 429344 125579
rect 429292 125536 429344 125545
rect 280804 125468 280856 125520
rect 281356 125468 281408 125520
rect 322296 124108 322348 124160
rect 579896 124108 579948 124160
rect 58440 122884 58492 122936
rect 60280 122884 60332 122936
rect 2780 122136 2832 122188
rect 6184 122136 6236 122188
rect 54668 120096 54720 120148
rect 59360 120096 59412 120148
rect 280804 120096 280856 120148
rect 281172 120096 281224 120148
rect 283840 120096 283892 120148
rect 491300 120096 491352 120148
rect 280896 118643 280948 118652
rect 280896 118609 280905 118643
rect 280905 118609 280939 118643
rect 280939 118609 280948 118643
rect 280896 118600 280948 118609
rect 56048 117308 56100 117360
rect 59360 117308 59412 117360
rect 283656 117308 283708 117360
rect 347872 117308 347924 117360
rect 7932 115991 7984 116000
rect 7932 115957 7941 115991
rect 7941 115957 7975 115991
rect 7975 115957 7984 115991
rect 7932 115948 7984 115957
rect 429292 115991 429344 116000
rect 429292 115957 429301 115991
rect 429301 115957 429335 115991
rect 429335 115957 429344 115991
rect 429292 115948 429344 115957
rect 280988 115880 281040 115932
rect 542360 115880 542412 115932
rect 542544 115880 542596 115932
rect 280804 113908 280856 113960
rect 281172 113908 281224 113960
rect 280804 112344 280856 112396
rect 281356 112344 281408 112396
rect 57152 111800 57204 111852
rect 59636 111800 59688 111852
rect 283748 111800 283800 111852
rect 433340 111800 433392 111852
rect 284024 109012 284076 109064
rect 423680 109012 423732 109064
rect 4068 107652 4120 107704
rect 55772 107652 55824 107704
rect 284024 107652 284076 107704
rect 411260 107652 411312 107704
rect 280804 106496 280856 106548
rect 281356 106496 281408 106548
rect 280896 106335 280948 106344
rect 280896 106301 280905 106335
rect 280905 106301 280939 106335
rect 280939 106301 280948 106335
rect 280896 106292 280948 106301
rect 284024 106292 284076 106344
rect 374092 106292 374144 106344
rect 8024 106267 8076 106276
rect 8024 106233 8033 106267
rect 8033 106233 8067 106267
rect 8067 106233 8076 106267
rect 8024 106224 8076 106233
rect 280804 106224 280856 106276
rect 281172 106224 281224 106276
rect 280896 106199 280948 106208
rect 280896 106165 280905 106199
rect 280905 106165 280939 106199
rect 280939 106165 280948 106199
rect 280896 106156 280948 106165
rect 6184 103504 6236 103556
rect 59360 103504 59412 103556
rect 283840 103504 283892 103556
rect 313280 103504 313332 103556
rect 299664 101439 299716 101448
rect 299664 101405 299673 101439
rect 299673 101405 299707 101439
rect 299707 101405 299716 101439
rect 299664 101396 299716 101405
rect 542636 101439 542688 101448
rect 542636 101405 542645 101439
rect 542645 101405 542679 101439
rect 542679 101405 542688 101439
rect 542636 101396 542688 101405
rect 55956 100716 56008 100768
rect 59360 100716 59412 100768
rect 284208 100716 284260 100768
rect 286232 100716 286284 100768
rect 283656 99356 283708 99408
rect 554044 99356 554096 99408
rect 8024 99331 8076 99340
rect 8024 99297 8033 99331
rect 8033 99297 8067 99331
rect 8067 99297 8076 99331
rect 8024 99288 8076 99297
rect 299664 99331 299716 99340
rect 299664 99297 299673 99331
rect 299673 99297 299707 99331
rect 299707 99297 299716 99331
rect 299664 99288 299716 99297
rect 542728 99288 542780 99340
rect 60096 98880 60148 98932
rect 62304 98880 62356 98932
rect 283840 97996 283892 98048
rect 409144 97996 409196 98048
rect 281080 96840 281132 96892
rect 280988 96636 281040 96688
rect 281080 96636 281132 96688
rect 429108 96568 429160 96620
rect 429384 96568 429436 96620
rect 280988 96543 281040 96552
rect 280988 96509 280997 96543
rect 280997 96509 281031 96543
rect 281031 96509 281040 96543
rect 280988 96500 281040 96509
rect 283840 95208 283892 95260
rect 389824 95208 389876 95260
rect 280804 94596 280856 94648
rect 281172 94596 281224 94648
rect 280804 94460 280856 94512
rect 281356 94460 281408 94512
rect 283840 93780 283892 93832
rect 290464 93780 290516 93832
rect 8116 90992 8168 91044
rect 59360 90992 59412 91044
rect 284024 89700 284076 89752
rect 469220 89700 469272 89752
rect 280988 89675 281040 89684
rect 280988 89641 280997 89675
rect 280997 89641 281031 89675
rect 281031 89641 281040 89675
rect 280988 89632 281040 89641
rect 283840 89632 283892 89684
rect 308496 89632 308548 89684
rect 501604 88272 501656 88324
rect 579896 88272 579948 88324
rect 283840 86980 283892 87032
rect 318064 86980 318116 87032
rect 280988 86912 281040 86964
rect 299664 86955 299716 86964
rect 299664 86921 299673 86955
rect 299673 86921 299707 86955
rect 299707 86921 299716 86955
rect 299664 86912 299716 86921
rect 287888 86232 287940 86284
rect 331312 86232 331364 86284
rect 283840 85552 283892 85604
rect 433432 85552 433484 85604
rect 280804 85008 280856 85060
rect 281448 85008 281500 85060
rect 280804 84872 280856 84924
rect 281356 84872 281408 84924
rect 283656 81404 283708 81456
rect 286508 81404 286560 81456
rect 429292 80044 429344 80096
rect 3976 79976 4028 80028
rect 55864 79976 55916 80028
rect 429384 79908 429436 79960
rect 284208 78684 284260 78736
rect 403624 78684 403676 78736
rect 10324 78616 10376 78668
rect 59360 78616 59412 78668
rect 280896 77299 280948 77308
rect 280896 77265 280905 77299
rect 280905 77265 280939 77299
rect 280939 77265 280948 77299
rect 280896 77256 280948 77265
rect 299664 77299 299716 77308
rect 299664 77265 299673 77299
rect 299673 77265 299707 77299
rect 299707 77265 299716 77299
rect 299664 77256 299716 77265
rect 62212 77231 62264 77240
rect 62212 77197 62221 77231
rect 62221 77197 62255 77231
rect 62255 77197 62264 77231
rect 62212 77188 62264 77197
rect 280988 77231 281040 77240
rect 280988 77197 280997 77231
rect 280997 77197 281031 77231
rect 281031 77197 281040 77231
rect 280988 77188 281040 77197
rect 294696 77188 294748 77240
rect 579620 77188 579672 77240
rect 280804 75284 280856 75336
rect 281356 75284 281408 75336
rect 280804 75148 280856 75200
rect 281448 75148 281500 75200
rect 55864 74536 55916 74588
rect 59360 74536 59412 74588
rect 284208 74536 284260 74588
rect 358820 74536 358872 74588
rect 284208 71748 284260 71800
rect 334624 71748 334676 71800
rect 280896 67668 280948 67720
rect 62304 67600 62356 67652
rect 283840 67600 283892 67652
rect 496084 67600 496136 67652
rect 280896 67575 280948 67584
rect 280896 67541 280905 67575
rect 280905 67541 280939 67575
rect 280939 67541 280948 67575
rect 280896 67532 280948 67541
rect 299664 67575 299716 67584
rect 299664 67541 299673 67575
rect 299673 67541 299707 67575
rect 299707 67541 299716 67575
rect 299664 67532 299716 67541
rect 542544 67532 542596 67584
rect 542728 67532 542780 67584
rect 280804 67396 280856 67448
rect 281448 67396 281500 67448
rect 280804 65424 280856 65476
rect 281356 65424 281408 65476
rect 55680 65288 55732 65340
rect 59360 65288 59412 65340
rect 407764 64812 407816 64864
rect 580172 64812 580224 64864
rect 283840 63520 283892 63572
rect 289912 63520 289964 63572
rect 283840 62024 283892 62076
rect 304356 62024 304408 62076
rect 299664 60979 299716 60988
rect 299664 60945 299673 60979
rect 299673 60945 299707 60979
rect 299707 60945 299716 60979
rect 299664 60936 299716 60945
rect 4804 60664 4856 60716
rect 59360 60664 59412 60716
rect 280988 60596 281040 60648
rect 429384 60596 429436 60648
rect 429568 60596 429620 60648
rect 283840 57944 283892 57996
rect 494704 57944 494756 57996
rect 281356 52708 281408 52760
rect 337384 51688 337436 51740
rect 538220 51688 538272 51740
rect 281448 51076 281500 51128
rect 280804 51008 280856 51060
rect 280988 51008 281040 51060
rect 281356 51008 281408 51060
rect 305644 50328 305696 50380
rect 459652 50328 459704 50380
rect 280896 48331 280948 48340
rect 280896 48297 280905 48331
rect 280905 48297 280939 48331
rect 280939 48297 280948 48331
rect 280896 48288 280948 48297
rect 280804 48220 280856 48272
rect 281356 48220 281408 48272
rect 318064 47540 318116 47592
rect 561680 47540 561732 47592
rect 283840 45568 283892 45620
rect 386420 45568 386472 45620
rect 287796 44820 287848 44872
rect 310520 44820 310572 44872
rect 62212 44276 62264 44328
rect 283840 44140 283892 44192
rect 506480 44140 506532 44192
rect 277032 43868 277084 43920
rect 60464 43800 60516 43852
rect 144184 43800 144236 43852
rect 61016 43732 61068 43784
rect 61292 43664 61344 43716
rect 187700 43664 187752 43716
rect 211068 43664 211120 43716
rect 283104 43664 283156 43716
rect 62028 43596 62080 43648
rect 223856 43596 223908 43648
rect 60004 43528 60056 43580
rect 227720 43528 227772 43580
rect 60280 43460 60332 43512
rect 333980 43460 334032 43512
rect 334624 43460 334676 43512
rect 534080 43460 534132 43512
rect 3424 43392 3476 43444
rect 57060 43392 57112 43444
rect 61476 43392 61528 43444
rect 362960 43392 363012 43444
rect 60372 42916 60424 42968
rect 64144 42916 64196 42968
rect 200028 42848 200080 42900
rect 286324 42848 286376 42900
rect 233516 42780 233568 42832
rect 429384 42780 429436 42832
rect 248420 42712 248472 42764
rect 286416 42712 286468 42764
rect 94228 42644 94280 42696
rect 285128 42644 285180 42696
rect 55772 42576 55824 42628
rect 160468 42576 160520 42628
rect 185124 42576 185176 42628
rect 290556 42576 290608 42628
rect 53104 42508 53156 42560
rect 146484 42508 146536 42560
rect 191012 42508 191064 42560
rect 291936 42508 291988 42560
rect 195060 42440 195112 42492
rect 287704 42440 287756 42492
rect 168288 42372 168340 42424
rect 286140 42372 286192 42424
rect 157248 42304 157300 42356
rect 286232 42304 286284 42356
rect 41328 42236 41380 42288
rect 96528 42236 96580 42288
rect 155868 42236 155920 42288
rect 287244 42236 287296 42288
rect 56232 42168 56284 42220
rect 154488 42168 154540 42220
rect 285956 42168 286008 42220
rect 56324 42100 56376 42152
rect 128452 42100 128504 42152
rect 286048 42100 286100 42152
rect 3516 42032 3568 42084
rect 88984 42032 89036 42084
rect 128360 42032 128412 42084
rect 580264 42032 580316 42084
rect 255412 41964 255464 42016
rect 285312 41964 285364 42016
rect 51724 41896 51776 41948
rect 258356 41896 258408 41948
rect 262128 41896 262180 41948
rect 288716 41896 288768 41948
rect 279424 41420 279476 41472
rect 284668 41420 284720 41472
rect 8944 41352 8996 41404
rect 88156 41352 88208 41404
rect 96528 41352 96580 41404
rect 216772 41352 216824 41404
rect 494704 41352 494756 41404
rect 580172 41352 580224 41404
rect 7564 41284 7616 41336
rect 127716 41284 127768 41336
rect 137008 41327 137060 41336
rect 137008 41293 137017 41327
rect 137017 41293 137051 41327
rect 137051 41293 137060 41327
rect 137008 41284 137060 41293
rect 270132 41284 270184 41336
rect 338120 41284 338172 41336
rect 88984 41216 89036 41268
rect 97172 41216 97224 41268
rect 106004 41216 106056 41268
rect 128360 41216 128412 41268
rect 181260 41216 181312 41268
rect 182088 41216 182140 41268
rect 57060 41148 57112 41200
rect 143540 41148 143592 41200
rect 198004 41148 198056 41200
rect 204904 41148 204956 41200
rect 11704 41080 11756 41132
rect 89260 41080 89312 41132
rect 103980 41080 104032 41132
rect 121460 41080 121512 41132
rect 158628 41080 158680 41132
rect 210884 41216 210936 41268
rect 229652 41216 229704 41268
rect 239404 41216 239456 41268
rect 257252 41216 257304 41268
rect 365720 41216 365772 41268
rect 208308 41148 208360 41200
rect 211804 41148 211856 41200
rect 239588 41148 239640 41200
rect 380900 41148 380952 41200
rect 234620 41080 234672 41132
rect 405740 41080 405792 41132
rect 3608 41012 3660 41064
rect 106924 41012 106976 41064
rect 139676 41012 139728 41064
rect 356060 41012 356112 41064
rect 128820 40944 128872 40996
rect 129648 40944 129700 40996
rect 153476 40944 153528 40996
rect 383660 40944 383712 40996
rect 2688 40876 2740 40928
rect 235540 40876 235592 40928
rect 245476 40876 245528 40928
rect 441620 40876 441672 40928
rect 87236 40808 87288 40860
rect 322940 40808 322992 40860
rect 83188 40740 83240 40792
rect 115204 40740 115256 40792
rect 164332 40740 164384 40792
rect 407764 40740 407816 40792
rect 111892 40672 111944 40724
rect 376760 40672 376812 40724
rect 240508 40196 240560 40248
rect 241244 40196 241296 40248
rect 249340 40128 249392 40180
rect 255964 40128 256016 40180
rect 63500 40060 63552 40112
rect 65524 40060 65576 40112
rect 69388 40060 69440 40112
rect 70308 40060 70360 40112
rect 70492 40060 70544 40112
rect 71688 40060 71740 40112
rect 84292 40060 84344 40112
rect 85488 40060 85540 40112
rect 91100 40060 91152 40112
rect 92296 40060 92348 40112
rect 110972 40060 111024 40112
rect 111708 40060 111760 40112
rect 114836 40060 114888 40112
rect 115848 40060 115900 40112
rect 118884 40060 118936 40112
rect 119896 40060 119948 40112
rect 125876 40060 125928 40112
rect 126796 40060 126848 40112
rect 129740 40060 129792 40112
rect 131028 40060 131080 40112
rect 132684 40060 132736 40112
rect 133788 40060 133840 40112
rect 135628 40060 135680 40112
rect 136456 40060 136508 40112
rect 136732 40060 136784 40112
rect 137928 40060 137980 40112
rect 142620 40060 142672 40112
rect 143448 40060 143500 40112
rect 149612 40060 149664 40112
rect 150348 40060 150400 40112
rect 157524 40060 157576 40112
rect 158536 40060 158588 40112
rect 163412 40060 163464 40112
rect 164148 40060 164200 40112
rect 167276 40060 167328 40112
rect 168196 40060 168248 40112
rect 170220 40060 170272 40112
rect 171048 40060 171100 40112
rect 171324 40060 171376 40112
rect 172336 40060 172388 40112
rect 174268 40060 174320 40112
rect 175188 40060 175240 40112
rect 178132 40060 178184 40112
rect 179236 40060 179288 40112
rect 182180 40060 182232 40112
rect 183376 40060 183428 40112
rect 189172 40060 189224 40112
rect 190368 40060 190420 40112
rect 195980 40060 196032 40112
rect 197176 40060 197228 40112
rect 202972 40060 203024 40112
rect 204076 40060 204128 40112
rect 209780 40060 209832 40112
rect 210976 40060 211028 40112
rect 212908 40060 212960 40112
rect 213736 40060 213788 40112
rect 215852 40060 215904 40112
rect 216588 40060 216640 40112
rect 220820 40060 220872 40112
rect 222108 40060 222160 40112
rect 230572 40060 230624 40112
rect 231768 40060 231820 40112
rect 243452 40060 243504 40112
rect 244188 40060 244240 40112
rect 244556 40060 244608 40112
rect 245476 40060 245528 40112
rect 254308 40060 254360 40112
rect 255228 40060 255280 40112
rect 269212 40060 269264 40112
rect 270408 40060 270460 40112
rect 279148 40060 279200 40112
rect 280068 40060 280120 40112
rect 95148 39992 95200 40044
rect 533344 39992 533396 40044
rect 14464 39924 14516 39976
rect 264244 39924 264296 39976
rect 265164 39924 265216 39976
rect 329104 39924 329156 39976
rect 81348 39856 81400 39908
rect 299756 39856 299808 39908
rect 82268 39788 82320 39840
rect 295984 39788 296036 39840
rect 74356 39720 74408 39772
rect 284944 39720 284996 39772
rect 219716 39652 219768 39704
rect 291844 39652 291896 39704
rect 60924 39380 60976 39432
rect 186320 39380 186372 39432
rect 263508 39380 263560 39432
rect 282000 39380 282052 39432
rect 59728 39312 59780 39364
rect 390652 39312 390704 39364
rect 135168 38632 135220 38684
rect 137008 38607 137060 38616
rect 137008 38573 137017 38607
rect 137017 38573 137051 38607
rect 137051 38573 137060 38607
rect 137008 38564 137060 38573
rect 135168 38496 135220 38548
rect 245568 38088 245620 38140
rect 283196 38156 283248 38208
rect 241428 38020 241480 38072
rect 281540 38088 281592 38140
rect 61384 37952 61436 38004
rect 193220 37952 193272 38004
rect 202788 37952 202840 38004
rect 281080 38020 281132 38072
rect 280988 37952 281040 38004
rect 339500 37952 339552 38004
rect 59636 37884 59688 37936
rect 425152 37884 425204 37936
rect 99012 37272 99064 37324
rect 99288 37272 99340 37324
rect 149060 37315 149112 37324
rect 149060 37281 149069 37315
rect 149069 37281 149103 37315
rect 149103 37281 149112 37315
rect 149060 37272 149112 37281
rect 179328 36660 179380 36712
rect 281448 36660 281500 36712
rect 58440 36592 58492 36644
rect 281540 36592 281592 36644
rect 60096 36524 60148 36576
rect 379520 36524 379572 36576
rect 280896 36456 280948 36508
rect 281356 36456 281408 36508
rect 3424 35844 3476 35896
rect 286508 35844 286560 35896
rect 58808 35300 58860 35352
rect 252560 35300 252612 35352
rect 263416 35300 263468 35352
rect 283748 35300 283800 35352
rect 58900 35232 58952 35284
rect 340880 35232 340932 35284
rect 62304 35164 62356 35216
rect 346400 35164 346452 35216
rect 62396 35096 62448 35148
rect 62396 34892 62448 34944
rect 219348 33872 219400 33924
rect 282368 33872 282420 33924
rect 59912 33804 59964 33856
rect 448520 33804 448572 33856
rect 146576 33779 146628 33788
rect 146576 33745 146585 33779
rect 146585 33745 146619 33779
rect 146619 33745 146628 33779
rect 146576 33736 146628 33745
rect 172336 33736 172388 33788
rect 572720 33736 572772 33788
rect 164148 33124 164200 33176
rect 168380 33124 168432 33176
rect 179144 32512 179196 32564
rect 270500 32512 270552 32564
rect 64788 32444 64840 32496
rect 223212 32444 223264 32496
rect 269028 32444 269080 32496
rect 280896 32444 280948 32496
rect 213736 32376 213788 32428
rect 483020 32376 483072 32428
rect 237656 31832 237708 31884
rect 237656 31696 237708 31748
rect 280068 31288 280120 31340
rect 287244 31288 287296 31340
rect 119896 31220 119948 31272
rect 307760 31220 307812 31272
rect 58532 31152 58584 31204
rect 295340 31152 295392 31204
rect 146208 31084 146260 31136
rect 226340 31084 226392 31136
rect 271788 31084 271840 31136
rect 546500 31084 546552 31136
rect 59084 31016 59136 31068
rect 438860 31016 438912 31068
rect 223212 30268 223264 30320
rect 580172 30268 580224 30320
rect 128268 29656 128320 29708
rect 276020 29656 276072 29708
rect 268936 29588 268988 29640
rect 563060 29588 563112 29640
rect 135168 28976 135220 29028
rect 137100 28976 137152 29028
rect 146668 28976 146720 29028
rect 231768 28568 231820 28620
rect 313372 28568 313424 28620
rect 124128 28500 124180 28552
rect 234620 28500 234672 28552
rect 153016 28432 153068 28484
rect 264980 28432 265032 28484
rect 60556 28364 60608 28416
rect 350540 28364 350592 28416
rect 141976 28296 142028 28348
rect 484400 28296 484452 28348
rect 158536 28228 158588 28280
rect 502432 28228 502484 28280
rect 99288 27548 99340 27600
rect 149060 27591 149112 27600
rect 149060 27557 149069 27591
rect 149069 27557 149103 27591
rect 149103 27557 149112 27591
rect 149060 27548 149112 27557
rect 150624 27548 150676 27600
rect 242164 27004 242216 27056
rect 283932 27004 283984 27056
rect 58716 26936 58768 26988
rect 245752 26936 245804 26988
rect 70308 26868 70360 26920
rect 558920 26868 558972 26920
rect 170956 25712 171008 25764
rect 282092 25712 282144 25764
rect 148968 25644 149020 25696
rect 281172 25644 281224 25696
rect 61200 25576 61252 25628
rect 236000 25576 236052 25628
rect 241244 25576 241296 25628
rect 500960 25576 501012 25628
rect 126796 25508 126848 25560
rect 391940 25508 391992 25560
rect 220728 24420 220780 24472
rect 283012 24420 283064 24472
rect 85488 24352 85540 24404
rect 233240 24352 233292 24404
rect 148876 24284 148928 24336
rect 318800 24284 318852 24336
rect 215208 24216 215260 24268
rect 401600 24216 401652 24268
rect 59176 24148 59228 24200
rect 280160 24148 280212 24200
rect 135076 24080 135128 24132
rect 467932 24080 467984 24132
rect 176568 22992 176620 23044
rect 283472 22992 283524 23044
rect 68928 22924 68980 22976
rect 248420 22924 248472 22976
rect 130936 22856 130988 22908
rect 336740 22856 336792 22908
rect 60832 22788 60884 22840
rect 324320 22788 324372 22840
rect 144828 22720 144880 22772
rect 466460 22720 466512 22772
rect 3148 22040 3200 22092
rect 146668 22040 146720 22092
rect 139216 21496 139268 21548
rect 252652 21496 252704 21548
rect 253848 21496 253900 21548
rect 320180 21496 320232 21548
rect 162676 21428 162728 21480
rect 282276 21428 282328 21480
rect 131028 21360 131080 21412
rect 546592 21360 546644 21412
rect 203984 20000 204036 20052
rect 280620 20000 280672 20052
rect 62396 19932 62448 19984
rect 162860 19932 162912 19984
rect 179236 19932 179288 19984
rect 516140 19932 516192 19984
rect 135168 19592 135220 19644
rect 135168 19320 135220 19372
rect 135168 19227 135220 19236
rect 135168 19193 135177 19227
rect 135177 19193 135211 19227
rect 135211 19193 135220 19227
rect 135168 19184 135220 19193
rect 129648 18844 129700 18896
rect 237564 18844 237616 18896
rect 143356 18776 143408 18828
rect 281632 18776 281684 18828
rect 182088 18708 182140 18760
rect 520372 18708 520424 18760
rect 175188 18640 175240 18692
rect 514760 18640 514812 18692
rect 58992 18572 59044 18624
rect 488540 18572 488592 18624
rect 149060 18003 149112 18012
rect 149060 17969 149069 18003
rect 149069 17969 149103 18003
rect 149103 17969 149112 18003
rect 149060 17960 149112 17969
rect 55956 17892 56008 17944
rect 579804 17892 579856 17944
rect 168196 17484 168248 17536
rect 269120 17484 269172 17536
rect 204076 17416 204128 17468
rect 532700 17416 532752 17468
rect 57520 17348 57572 17400
rect 443092 17348 443144 17400
rect 111708 17280 111760 17332
rect 505100 17280 505152 17332
rect 103428 17212 103480 17264
rect 513380 17212 513432 17264
rect 231768 16124 231820 16176
rect 283564 16124 283616 16176
rect 118608 16056 118660 16108
rect 247132 16056 247184 16108
rect 270408 16056 270460 16108
rect 291200 16056 291252 16108
rect 304264 16056 304316 16108
rect 528652 16056 528704 16108
rect 59268 15988 59320 16040
rect 309140 15988 309192 16040
rect 115848 15920 115900 15972
rect 414020 15920 414072 15972
rect 197176 15852 197228 15904
rect 510620 15852 510672 15904
rect 210976 14628 211028 14680
rect 321560 14628 321612 14680
rect 71596 14560 71648 14612
rect 236092 14560 236144 14612
rect 240048 14560 240100 14612
rect 281264 14560 281316 14612
rect 140688 14492 140740 14544
rect 371240 14492 371292 14544
rect 121368 14424 121420 14476
rect 569960 14424 570012 14476
rect 182088 13744 182140 13796
rect 185124 13744 185176 13796
rect 256516 13200 256568 13252
rect 283380 13200 283432 13252
rect 190368 13132 190420 13184
rect 343640 13132 343692 13184
rect 137928 13064 137980 13116
rect 553400 13064 553452 13116
rect 554044 13064 554096 13116
rect 560300 13064 560352 13116
rect 149060 12452 149112 12504
rect 237472 12452 237524 12504
rect 237748 12452 237800 12504
rect 149244 12248 149296 12300
rect 166908 12044 166960 12096
rect 247040 12044 247092 12096
rect 136456 11976 136508 12028
rect 167000 11976 167052 12028
rect 183376 11976 183428 12028
rect 283012 11976 283064 12028
rect 131396 11908 131448 11960
rect 281908 11908 281960 11960
rect 133604 11840 133656 11892
rect 237472 11840 237524 11892
rect 252468 11840 252520 11892
rect 408592 11840 408644 11892
rect 60740 11772 60792 11824
rect 299480 11772 299532 11824
rect 308404 11772 308456 11824
rect 507860 11772 507912 11824
rect 58624 11704 58676 11756
rect 444380 11704 444432 11756
rect 150716 11679 150768 11688
rect 150716 11645 150725 11679
rect 150725 11645 150759 11679
rect 150759 11645 150768 11679
rect 150716 11636 150768 11645
rect 385684 10956 385736 11008
rect 389180 10956 389232 11008
rect 409144 10956 409196 11008
rect 409880 10956 409932 11008
rect 205548 10684 205600 10736
rect 335360 10684 335412 10736
rect 172428 10616 172480 10668
rect 342260 10616 342312 10668
rect 193128 10548 193180 10600
rect 364340 10548 364392 10600
rect 171048 10480 171100 10532
rect 353300 10480 353352 10532
rect 155776 10412 155828 10464
rect 349160 10412 349212 10464
rect 371884 10412 371936 10464
rect 385040 10412 385092 10464
rect 92296 10344 92348 10396
rect 356152 10344 356204 10396
rect 364984 10344 365036 10396
rect 382280 10344 382332 10396
rect 389824 10344 389876 10396
rect 407120 10344 407172 10396
rect 60648 10276 60700 10328
rect 328460 10276 328512 10328
rect 356704 10276 356756 10328
rect 463700 10276 463752 10328
rect 99196 9707 99248 9716
rect 99196 9673 99205 9707
rect 99205 9673 99239 9707
rect 99239 9673 99248 9707
rect 99196 9664 99248 9673
rect 134892 9664 134944 9716
rect 234528 9664 234580 9716
rect 234804 9664 234856 9716
rect 169668 9596 169720 9648
rect 250352 9596 250404 9648
rect 257436 9596 257488 9648
rect 288624 9596 288676 9648
rect 162768 9528 162820 9580
rect 243176 9528 243228 9580
rect 245476 9528 245528 9580
rect 303804 9528 303856 9580
rect 187608 9460 187660 9512
rect 318064 9460 318116 9512
rect 122748 9392 122800 9444
rect 275284 9392 275336 9444
rect 113088 9324 113140 9376
rect 321652 9324 321704 9376
rect 53380 9256 53432 9308
rect 278872 9256 278924 9308
rect 180708 9188 180760 9240
rect 225328 9188 225380 9240
rect 239404 9188 239456 9240
rect 478696 9188 478748 9240
rect 53196 9120 53248 9172
rect 294328 9120 294380 9172
rect 54668 9052 54720 9104
rect 315764 9052 315816 9104
rect 322204 9052 322256 9104
rect 360936 9052 360988 9104
rect 53288 8984 53340 9036
rect 326436 8984 326488 9036
rect 126888 8916 126940 8968
rect 228916 8916 228968 8968
rect 256608 8916 256660 8968
rect 575020 8916 575072 8968
rect 196808 8848 196860 8900
rect 251180 8848 251232 8900
rect 264612 8848 264664 8900
rect 289820 8848 289872 8900
rect 189632 8780 189684 8832
rect 241520 8780 241572 8832
rect 218152 8712 218204 8764
rect 237380 8712 237432 8764
rect 208216 7964 208268 8016
rect 214656 7964 214708 8016
rect 159916 7896 159968 7948
rect 282920 7896 282972 7948
rect 184848 7828 184900 7880
rect 395436 7828 395488 7880
rect 61108 7760 61160 7812
rect 221740 7760 221792 7812
rect 224868 7760 224920 7812
rect 545304 7760 545356 7812
rect 213828 7692 213880 7744
rect 538128 7692 538180 7744
rect 65524 7624 65576 7676
rect 399024 7624 399076 7676
rect 204168 7556 204220 7608
rect 555976 7556 556028 7608
rect 2964 7352 3016 7404
rect 6184 7352 6236 7404
rect 212264 6808 212316 6860
rect 284576 6808 284628 6860
rect 192024 6740 192076 6792
rect 281816 6740 281868 6792
rect 144460 6672 144512 6724
rect 223672 6672 223724 6724
rect 251088 6672 251140 6724
rect 388260 6672 388312 6724
rect 53656 6604 53708 6656
rect 177764 6604 177816 6656
rect 182548 6604 182600 6656
rect 245660 6604 245712 6656
rect 266176 6604 266228 6656
rect 404912 6604 404964 6656
rect 54852 6536 54904 6588
rect 272892 6536 272944 6588
rect 274548 6536 274600 6588
rect 365812 6536 365864 6588
rect 55680 6468 55732 6520
rect 279976 6468 280028 6520
rect 53748 6400 53800 6452
rect 195612 6400 195664 6452
rect 226248 6400 226300 6452
rect 495348 6400 495400 6452
rect 133788 6332 133840 6384
rect 422760 6332 422812 6384
rect 92388 6264 92440 6316
rect 383568 6264 383620 6316
rect 54944 6196 54996 6248
rect 213460 6196 213512 6248
rect 241336 6196 241388 6248
rect 541716 6196 541768 6248
rect 119988 6128 120040 6180
rect 440608 6128 440660 6180
rect 244188 6060 244240 6112
rect 306196 6060 306248 6112
rect 267004 5992 267056 6044
rect 284392 5992 284444 6044
rect 277676 5924 277728 5976
rect 288532 5924 288584 5976
rect 180156 5176 180208 5228
rect 198740 5176 198792 5228
rect 183468 5108 183520 5160
rect 215852 5108 215904 5160
rect 222108 5108 222160 5160
rect 230112 5108 230164 5160
rect 241980 5108 242032 5160
rect 283656 5108 283708 5160
rect 132408 5040 132460 5092
rect 201500 5040 201552 5092
rect 208676 5040 208728 5092
rect 260840 5040 260892 5092
rect 267648 5040 267700 5092
rect 271696 5040 271748 5092
rect 143448 4972 143500 5024
rect 274088 4972 274140 5024
rect 278688 4972 278740 5024
rect 551192 4972 551244 5024
rect 197268 4904 197320 4956
rect 523868 4904 523920 4956
rect 108948 4836 109000 4888
rect 453672 4836 453724 4888
rect 71688 4768 71740 4820
rect 579804 4768 579856 4820
rect 281540 4156 281592 4208
rect 282460 4156 282512 4208
rect 55036 4088 55088 4140
rect 161112 4088 161164 4140
rect 239588 4088 239640 4140
rect 240048 4088 240100 4140
rect 255044 4088 255096 4140
rect 287152 4088 287204 4140
rect 514024 4088 514076 4140
rect 514576 4088 514628 4140
rect 57796 4020 57848 4072
rect 164700 4020 164752 4072
rect 205088 4020 205140 4072
rect 279424 4020 279476 4072
rect 281540 4020 281592 4072
rect 282184 4020 282236 4072
rect 403624 4020 403676 4072
rect 56416 3952 56468 4004
rect 176476 3952 176528 4004
rect 183744 3952 183796 4004
rect 285772 3952 285824 4004
rect 407764 3952 407816 4004
rect 435824 3952 435876 4004
rect 57888 3884 57940 3936
rect 186044 3884 186096 3936
rect 199200 3884 199252 3936
rect 281724 3884 281776 3936
rect 356152 3884 356204 3936
rect 357348 3884 357400 3936
rect 390652 3884 390704 3936
rect 391848 3884 391900 3936
rect 408500 3884 408552 3936
rect 409696 3884 409748 3936
rect 432328 3884 432380 3936
rect 57152 3816 57204 3868
rect 190828 3816 190880 3868
rect 217048 3816 217100 3868
rect 242164 3816 242216 3868
rect 255964 3816 256016 3868
rect 417976 3816 418028 3868
rect 57612 3748 57664 3800
rect 222936 3748 222988 3800
rect 255228 3748 255280 3800
rect 421564 3748 421616 3800
rect 53564 3680 53616 3732
rect 244372 3680 244424 3732
rect 251456 3680 251508 3732
rect 284484 3680 284536 3732
rect 285220 3680 285272 3732
rect 475108 3680 475160 3732
rect 502984 3680 503036 3732
rect 57704 3612 57756 3664
rect 198004 3612 198056 3664
rect 204904 3612 204956 3664
rect 425060 3612 425112 3664
rect 459652 3612 459704 3664
rect 460848 3612 460900 3664
rect 467104 3612 467156 3664
rect 497740 3612 497792 3664
rect 64144 3544 64196 3596
rect 206284 3544 206336 3596
rect 216588 3544 216640 3596
rect 471520 3544 471572 3596
rect 496084 3544 496136 3596
rect 502340 3544 502392 3596
rect 502432 3544 502484 3596
rect 503628 3544 503680 3596
rect 520280 3612 520332 3664
rect 521476 3612 521528 3664
rect 528652 3612 528704 3664
rect 529848 3612 529900 3664
rect 552388 3544 552440 3596
rect 563152 3544 563204 3596
rect 564348 3544 564400 3596
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 55128 3408 55180 3460
rect 62488 3340 62540 3392
rect 115204 3476 115256 3528
rect 425152 3476 425204 3528
rect 426348 3476 426400 3528
rect 433340 3476 433392 3528
rect 434628 3476 434680 3528
rect 435364 3476 435416 3528
rect 567844 3476 567896 3528
rect 574744 3476 574796 3528
rect 581000 3476 581052 3528
rect 128452 3408 128504 3460
rect 129004 3408 129056 3460
rect 136088 3408 136140 3460
rect 136548 3408 136600 3460
rect 136732 3408 136784 3460
rect 137284 3408 137336 3460
rect 138480 3408 138532 3460
rect 139308 3408 139360 3460
rect 140872 3408 140924 3460
rect 142068 3408 142120 3460
rect 144184 3408 144236 3460
rect 145656 3408 145708 3460
rect 148048 3408 148100 3460
rect 148968 3408 149020 3460
rect 150716 3408 150768 3460
rect 151544 3408 151596 3460
rect 153936 3408 153988 3460
rect 154488 3408 154540 3460
rect 155132 3408 155184 3460
rect 155868 3408 155920 3460
rect 122748 3340 122800 3392
rect 56508 3272 56560 3324
rect 127808 3272 127860 3324
rect 128268 3272 128320 3324
rect 150348 3340 150400 3392
rect 482284 3408 482336 3460
rect 482376 3408 482428 3460
rect 496544 3408 496596 3460
rect 497464 3408 497516 3460
rect 509608 3408 509660 3460
rect 514576 3408 514628 3460
rect 577412 3408 577464 3460
rect 156328 3340 156380 3392
rect 157248 3340 157300 3392
rect 157524 3340 157576 3392
rect 158628 3340 158680 3392
rect 158720 3340 158772 3392
rect 160008 3340 160060 3392
rect 175372 3340 175424 3392
rect 176568 3340 176620 3392
rect 181352 3340 181404 3392
rect 182088 3340 182140 3392
rect 183560 3340 183612 3392
rect 184848 3340 184900 3392
rect 231308 3340 231360 3392
rect 231768 3340 231820 3392
rect 252560 3340 252612 3392
rect 253848 3340 253900 3392
rect 261024 3340 261076 3392
rect 262128 3340 262180 3392
rect 262220 3340 262272 3392
rect 263508 3340 263560 3392
rect 285680 3340 285732 3392
rect 287060 3340 287112 3392
rect 288348 3340 288400 3392
rect 296720 3340 296772 3392
rect 297916 3340 297968 3392
rect 313280 3340 313332 3392
rect 314568 3340 314620 3392
rect 321560 3340 321612 3392
rect 322848 3340 322900 3392
rect 347780 3340 347832 3392
rect 349068 3340 349120 3392
rect 365720 3340 365772 3392
rect 366916 3340 366968 3392
rect 374000 3340 374052 3392
rect 375196 3340 375248 3392
rect 428740 3340 428792 3392
rect 443000 3340 443052 3392
rect 444196 3340 444248 3392
rect 467932 3340 467984 3392
rect 469128 3340 469180 3392
rect 150440 3272 150492 3324
rect 240784 3272 240836 3324
rect 241428 3272 241480 3324
rect 259828 3272 259880 3324
rect 285864 3272 285916 3324
rect 142068 3204 142120 3256
rect 268108 3204 268160 3256
rect 269028 3204 269080 3256
rect 276480 3204 276532 3256
rect 281540 3204 281592 3256
rect 130200 3136 130252 3188
rect 258632 3136 258684 3188
rect 99196 3000 99248 3052
rect 122748 3000 122800 3052
rect 132592 3000 132644 3052
rect 207480 3000 207532 3052
rect 208308 3000 208360 3052
rect 165896 2932 165948 2984
rect 166908 2932 166960 2984
rect 193220 2864 193272 2916
rect 194416 2864 194468 2916
rect 153108 2796 153160 2848
rect 194508 2796 194560 2848
rect 280068 2796 280120 2848
rect 490564 2796 490616 2848
rect 193220 2728 193272 2780
rect 152740 595 152792 604
rect 152740 561 152749 595
rect 152749 561 152783 595
rect 152783 561 152792 595
rect 152740 552 152792 561
rect 186320 552 186372 604
rect 187240 552 187292 604
rect 187700 552 187752 604
rect 188436 552 188488 604
rect 236092 552 236144 604
rect 237196 552 237248 604
rect 237564 552 237616 604
rect 238392 552 238444 604
rect 280160 552 280212 604
rect 281264 552 281316 604
rect 316040 552 316092 604
rect 316960 552 317012 604
rect 318800 552 318852 604
rect 319260 552 319312 604
rect 322940 552 322992 604
rect 324044 552 324096 604
rect 324320 552 324372 604
rect 325240 552 325292 604
rect 393320 552 393372 604
rect 394240 552 394292 604
rect 396080 552 396132 604
rect 396632 552 396684 604
rect 401600 552 401652 604
rect 402520 552 402572 604
rect 412640 552 412692 604
rect 413284 552 413336 604
rect 415400 552 415452 604
rect 415676 552 415728 604
rect 418160 552 418212 604
rect 419172 552 419224 604
rect 419540 552 419592 604
rect 420368 552 420420 604
rect 547880 552 547932 604
rect 548892 552 548944 604
rect 549260 552 549312 604
rect 550088 552 550140 604
rect 556160 552 556212 604
rect 557172 552 557224 604
rect 581092 552 581144 604
rect 582196 552 582248 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 700398 24348 703520
rect 40512 700466 40540 703520
rect 72988 700534 73016 703520
rect 72976 700528 73028 700534
rect 72976 700470 73028 700476
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3330 682272 3386 682281
rect 3330 682207 3386 682216
rect 3344 681766 3372 682207
rect 3332 681760 3384 681766
rect 3332 681702 3384 681708
rect 4804 681760 4856 681766
rect 4804 681702 4856 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3330 653576 3386 653585
rect 3330 653511 3386 653520
rect 3344 652905 3372 653511
rect 3330 652896 3386 652905
rect 3330 652831 3386 652840
rect 4066 624880 4122 624889
rect 4066 624815 4122 624824
rect 4080 623830 4108 624815
rect 4068 623824 4120 623830
rect 4068 623766 4120 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 4066 567352 4122 567361
rect 4066 567287 4122 567296
rect 4080 567254 4108 567287
rect 4068 567248 4120 567254
rect 4068 567190 4120 567196
rect 4066 553072 4122 553081
rect 4066 553007 4122 553016
rect 4080 552090 4108 553007
rect 4068 552084 4120 552090
rect 4068 552026 4120 552032
rect 3974 538656 4030 538665
rect 3974 538591 4030 538600
rect 3988 538490 4016 538591
rect 3976 538484 4028 538490
rect 3976 538426 4028 538432
rect 3882 509960 3938 509969
rect 3882 509895 3938 509904
rect 3896 509318 3924 509895
rect 3884 509312 3936 509318
rect 3884 509254 3936 509260
rect 4066 495544 4122 495553
rect 4066 495479 4068 495488
rect 4120 495479 4122 495488
rect 4068 495450 4120 495456
rect 3330 481128 3386 481137
rect 3330 481063 3386 481072
rect 3344 480622 3372 481063
rect 3332 480616 3384 480622
rect 3332 480558 3384 480564
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 3146 294400 3202 294409
rect 3146 294335 3202 294344
rect 3160 294030 3188 294335
rect 3148 294024 3200 294030
rect 3148 293966 3200 293972
rect 1308 261452 1360 261458
rect 1308 261394 1360 261400
rect 1320 3534 1348 261394
rect 2964 223508 3016 223514
rect 2964 223450 3016 223456
rect 2976 222601 3004 223450
rect 2962 222592 3018 222601
rect 2962 222527 3018 222536
rect 3332 165572 3384 165578
rect 3332 165514 3384 165520
rect 3344 165073 3372 165514
rect 3330 165064 3386 165073
rect 3330 164999 3386 165008
rect 2780 122188 2832 122194
rect 2780 122130 2832 122136
rect 2792 122097 2820 122130
rect 2778 122088 2834 122097
rect 2778 122023 2834 122032
rect 3436 43450 3464 452367
rect 3790 438016 3846 438025
rect 3790 437951 3846 437960
rect 3804 437510 3832 437951
rect 3792 437504 3844 437510
rect 3792 437446 3844 437452
rect 4066 423736 4122 423745
rect 4066 423671 4068 423680
rect 4120 423671 4122 423680
rect 4068 423642 4120 423648
rect 4066 395040 4122 395049
rect 4066 394975 4122 394984
rect 4080 394738 4108 394975
rect 4068 394732 4120 394738
rect 4068 394674 4120 394680
rect 3974 380624 4030 380633
rect 3974 380559 4030 380568
rect 3988 379574 4016 380559
rect 3976 379568 4028 379574
rect 3976 379510 4028 379516
rect 4066 366208 4122 366217
rect 4066 366143 4122 366152
rect 4080 365770 4108 366143
rect 4068 365764 4120 365770
rect 4068 365706 4120 365712
rect 4066 337512 4122 337521
rect 4066 337447 4122 337456
rect 4080 336802 4108 337447
rect 4068 336796 4120 336802
rect 4068 336738 4120 336744
rect 3606 323096 3662 323105
rect 3606 323031 3662 323040
rect 3516 265736 3568 265742
rect 3516 265678 3568 265684
rect 3528 64569 3556 265678
rect 3620 223582 3648 323031
rect 4066 308816 4122 308825
rect 4066 308751 4122 308760
rect 4080 307834 4108 308751
rect 4068 307828 4120 307834
rect 4068 307770 4120 307776
rect 3698 280120 3754 280129
rect 3698 280055 3754 280064
rect 3608 223576 3660 223582
rect 3608 223518 3660 223524
rect 3712 189038 3740 280055
rect 3884 266348 3936 266354
rect 3884 266290 3936 266296
rect 3896 265713 3924 266290
rect 3882 265704 3938 265713
rect 3882 265639 3938 265648
rect 4066 251288 4122 251297
rect 4066 251223 4068 251232
rect 4120 251223 4122 251232
rect 4068 251194 4120 251200
rect 4068 237380 4120 237386
rect 4068 237322 4120 237328
rect 4080 237017 4108 237322
rect 4066 237008 4122 237017
rect 4066 236943 4122 236952
rect 3700 189032 3752 189038
rect 3700 188974 3752 188980
rect 4066 180704 4122 180713
rect 4066 180639 4122 180648
rect 4080 179489 4108 180639
rect 4066 179480 4122 179489
rect 4066 179415 4122 179424
rect 3606 150784 3662 150793
rect 3606 150719 3662 150728
rect 3514 64560 3570 64569
rect 3514 64495 3570 64504
rect 3514 50144 3570 50153
rect 3514 50079 3570 50088
rect 3424 43444 3476 43450
rect 3424 43386 3476 43392
rect 3528 42090 3556 50079
rect 3516 42084 3568 42090
rect 3516 42026 3568 42032
rect 3620 41070 3648 150719
rect 3974 136368 4030 136377
rect 3974 136303 4030 136312
rect 3988 135318 4016 136303
rect 3976 135312 4028 135318
rect 3976 135254 4028 135260
rect 4068 107704 4120 107710
rect 4066 107672 4068 107681
rect 4120 107672 4122 107681
rect 4066 107607 4122 107616
rect 3976 80028 4028 80034
rect 3976 79970 4028 79976
rect 3988 78985 4016 79970
rect 3974 78976 4030 78985
rect 3974 78911 4030 78920
rect 4816 60722 4844 681702
rect 8128 679046 8156 685850
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654158 8064 663734
rect 8024 654152 8076 654158
rect 8024 654094 8076 654100
rect 8208 654152 8260 654158
rect 8208 654094 8260 654100
rect 8220 644450 8248 654094
rect 8036 644422 8248 644450
rect 8036 634846 8064 644422
rect 8024 634840 8076 634846
rect 8024 634782 8076 634788
rect 8208 634840 8260 634846
rect 8208 634782 8260 634788
rect 8220 625138 8248 634782
rect 8036 625110 8248 625138
rect 6184 623824 6236 623830
rect 6184 623766 6236 623772
rect 6196 260846 6224 623766
rect 8036 615534 8064 625110
rect 8024 615528 8076 615534
rect 8024 615470 8076 615476
rect 8208 615528 8260 615534
rect 8208 615470 8260 615476
rect 8220 605826 8248 615470
rect 14556 610020 14608 610026
rect 14556 609962 14608 609968
rect 8036 605798 8248 605826
rect 8036 596222 8064 605798
rect 8024 596216 8076 596222
rect 8208 596216 8260 596222
rect 8024 596158 8076 596164
rect 8128 596164 8208 596170
rect 8128 596158 8260 596164
rect 8128 596142 8248 596158
rect 8128 591954 8156 596142
rect 8036 591926 8156 591954
rect 8036 589286 8064 591926
rect 8024 589280 8076 589286
rect 8024 589222 8076 589228
rect 8024 579760 8076 579766
rect 7944 579708 8024 579714
rect 7944 579702 8076 579708
rect 7944 579686 8064 579702
rect 7944 579630 7972 579686
rect 7932 579624 7984 579630
rect 7932 579566 7984 579572
rect 8116 579624 8168 579630
rect 8116 579566 8168 579572
rect 8128 562970 8156 579566
rect 7932 562964 7984 562970
rect 7932 562906 7984 562912
rect 8116 562964 8168 562970
rect 8116 562906 8168 562912
rect 7944 553330 7972 562906
rect 7944 553302 8064 553330
rect 8036 550594 8064 553302
rect 8024 550588 8076 550594
rect 8024 550530 8076 550536
rect 8208 541000 8260 541006
rect 8208 540942 8260 540948
rect 8220 534018 8248 540942
rect 10324 538484 10376 538490
rect 10324 538426 10376 538432
rect 8128 533990 8248 534018
rect 8128 531321 8156 533990
rect 8114 531312 8170 531321
rect 8114 531247 8170 531256
rect 8390 531312 8446 531321
rect 8390 531247 8446 531256
rect 8404 521694 8432 531247
rect 8208 521688 8260 521694
rect 8208 521630 8260 521636
rect 8392 521688 8444 521694
rect 8392 521630 8444 521636
rect 8220 514706 8248 521630
rect 8128 514678 8248 514706
rect 8128 512009 8156 514678
rect 8114 512000 8170 512009
rect 8114 511935 8170 511944
rect 8390 512000 8446 512009
rect 8390 511935 8446 511944
rect 8404 502382 8432 511935
rect 8208 502376 8260 502382
rect 8208 502318 8260 502324
rect 8392 502376 8444 502382
rect 8392 502318 8444 502324
rect 8220 495394 8248 502318
rect 8128 495366 8248 495394
rect 8128 492658 8156 495366
rect 7932 492652 7984 492658
rect 7932 492594 7984 492600
rect 8116 492652 8168 492658
rect 8116 492594 8168 492600
rect 7944 483041 7972 492594
rect 7930 483032 7986 483041
rect 7930 482967 7986 482976
rect 8206 483032 8262 483041
rect 8206 482967 8262 482976
rect 8220 476082 8248 482967
rect 8036 476054 8248 476082
rect 8036 473346 8064 476054
rect 8024 473340 8076 473346
rect 8024 473282 8076 473288
rect 8116 473340 8168 473346
rect 8116 473282 8168 473288
rect 8128 463706 8156 473282
rect 8128 463678 8248 463706
rect 8220 456770 8248 463678
rect 8036 456742 8248 456770
rect 8036 447166 8064 456742
rect 8024 447160 8076 447166
rect 8024 447102 8076 447108
rect 8116 447092 8168 447098
rect 8116 447034 8168 447040
rect 8128 444378 8156 447034
rect 7840 444372 7892 444378
rect 7840 444314 7892 444320
rect 8116 444372 8168 444378
rect 8116 444314 8168 444320
rect 7852 434761 7880 444314
rect 7838 434752 7894 434761
rect 7838 434687 7894 434696
rect 8022 434752 8078 434761
rect 8022 434687 8078 434696
rect 8036 427922 8064 434687
rect 8024 427916 8076 427922
rect 8024 427858 8076 427864
rect 8024 427780 8076 427786
rect 8024 427722 8076 427728
rect 8036 418198 8064 427722
rect 8024 418192 8076 418198
rect 8024 418134 8076 418140
rect 8208 418192 8260 418198
rect 8208 418134 8260 418140
rect 8220 408490 8248 418134
rect 8036 408462 8248 408490
rect 8036 398954 8064 408462
rect 8024 398948 8076 398954
rect 8024 398890 8076 398896
rect 8036 390590 8064 390621
rect 8024 390584 8076 390590
rect 7852 390532 8024 390538
rect 7852 390526 8076 390532
rect 7852 390510 8064 390526
rect 7852 380934 7880 390510
rect 7840 380928 7892 380934
rect 7840 380870 7892 380876
rect 8024 380928 8076 380934
rect 8024 380870 8076 380876
rect 8036 369918 8064 380870
rect 8024 369912 8076 369918
rect 8024 369854 8076 369860
rect 7932 369844 7984 369850
rect 7932 369786 7984 369792
rect 7944 360194 7972 369786
rect 7932 360188 7984 360194
rect 7932 360130 7984 360136
rect 8116 360188 8168 360194
rect 8116 360130 8168 360136
rect 8128 357406 8156 360130
rect 8116 357400 8168 357406
rect 8116 357342 8168 357348
rect 8024 347812 8076 347818
rect 8024 347754 8076 347760
rect 8036 341018 8064 347754
rect 8024 341012 8076 341018
rect 8024 340954 8076 340960
rect 8024 336864 8076 336870
rect 8024 336806 8076 336812
rect 8036 336666 8064 336806
rect 8024 336660 8076 336666
rect 8024 336602 8076 336608
rect 7932 327140 7984 327146
rect 7932 327082 7984 327088
rect 7944 321502 7972 327082
rect 7932 321496 7984 321502
rect 7932 321438 7984 321444
rect 8208 321496 8260 321502
rect 8208 321438 8260 321444
rect 8220 309262 8248 321438
rect 7932 309256 7984 309262
rect 8208 309256 8260 309262
rect 7984 309204 8064 309210
rect 7932 309198 8064 309204
rect 8208 309198 8260 309204
rect 7944 309182 8064 309198
rect 8036 302326 8064 309182
rect 8024 302320 8076 302326
rect 8024 302262 8076 302268
rect 8116 302116 8168 302122
rect 8116 302058 8168 302064
rect 7564 294024 7616 294030
rect 7564 293966 7616 293972
rect 6276 268116 6328 268122
rect 6276 268058 6328 268064
rect 6184 260840 6236 260846
rect 6184 260782 6236 260788
rect 4894 194576 4950 194585
rect 4894 194511 4950 194520
rect 4908 193905 4936 194511
rect 4894 193896 4950 193905
rect 4894 193831 4950 193840
rect 6288 165578 6316 268058
rect 6276 165572 6328 165578
rect 6276 165514 6328 165520
rect 6184 150476 6236 150482
rect 6184 150418 6236 150424
rect 6196 122194 6224 150418
rect 6184 122188 6236 122194
rect 6184 122130 6236 122136
rect 6184 103556 6236 103562
rect 6184 103498 6236 103504
rect 4804 60716 4856 60722
rect 4804 60658 4856 60664
rect 3608 41064 3660 41070
rect 3608 41006 3660 41012
rect 2688 40928 2740 40934
rect 2688 40870 2740 40876
rect 2700 3534 2728 40870
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 6196 7410 6224 103498
rect 7576 41342 7604 293966
rect 8128 292618 8156 302058
rect 8128 292590 8248 292618
rect 8220 289814 8248 292590
rect 8208 289808 8260 289814
rect 8208 289750 8260 289756
rect 8116 280220 8168 280226
rect 8116 280162 8168 280168
rect 8128 273358 8156 280162
rect 8116 273352 8168 273358
rect 8116 273294 8168 273300
rect 8116 273148 8168 273154
rect 8116 273090 8168 273096
rect 8128 244202 8156 273090
rect 8944 251252 8996 251258
rect 8944 251194 8996 251200
rect 8036 244174 8156 244202
rect 8036 231878 8064 244174
rect 7932 231872 7984 231878
rect 7932 231814 7984 231820
rect 8024 231872 8076 231878
rect 8024 231814 8076 231820
rect 7944 224890 7972 231814
rect 7944 224862 8064 224890
rect 8036 222154 8064 224862
rect 8024 222148 8076 222154
rect 8024 222090 8076 222096
rect 8116 215212 8168 215218
rect 8116 215154 8168 215160
rect 8128 205766 8156 215154
rect 8116 205760 8168 205766
rect 8116 205702 8168 205708
rect 7932 205624 7984 205630
rect 7932 205566 7984 205572
rect 7944 201482 7972 205566
rect 7932 201476 7984 201482
rect 7932 201418 7984 201424
rect 7932 193180 7984 193186
rect 7932 193122 7984 193128
rect 7944 191842 7972 193122
rect 7944 191814 8064 191842
rect 8036 186386 8064 191814
rect 8024 186380 8076 186386
rect 8024 186322 8076 186328
rect 8116 186244 8168 186250
rect 8116 186186 8168 186192
rect 8128 176798 8156 186186
rect 8116 176792 8168 176798
rect 8116 176734 8168 176740
rect 8024 176588 8076 176594
rect 8024 176530 8076 176536
rect 8036 164218 8064 176530
rect 8024 164212 8076 164218
rect 8024 164154 8076 164160
rect 8116 164212 8168 164218
rect 8116 164154 8168 164160
rect 8128 154578 8156 164154
rect 8128 154550 8248 154578
rect 8220 147642 8248 154550
rect 8036 147614 8248 147642
rect 8036 144906 8064 147614
rect 8024 144900 8076 144906
rect 8024 144842 8076 144848
rect 8116 144900 8168 144906
rect 8116 144842 8168 144848
rect 8128 135266 8156 144842
rect 8128 135238 8248 135266
rect 8220 128330 8248 135238
rect 8036 128302 8248 128330
rect 8036 125594 8064 128302
rect 8024 125588 8076 125594
rect 8024 125530 8076 125536
rect 7932 116000 7984 116006
rect 7932 115942 7984 115948
rect 7944 109018 7972 115942
rect 7944 108990 8064 109018
rect 8036 106282 8064 108990
rect 8024 106276 8076 106282
rect 8024 106218 8076 106224
rect 8024 99340 8076 99346
rect 8024 99282 8076 99288
rect 8036 96642 8064 99282
rect 8036 96614 8156 96642
rect 8128 91050 8156 96614
rect 8116 91044 8168 91050
rect 8116 90986 8168 90992
rect 8956 41410 8984 251194
rect 10336 78674 10364 538426
rect 11704 480616 11756 480622
rect 11704 480558 11756 480564
rect 10324 78668 10376 78674
rect 10324 78610 10376 78616
rect 8944 41404 8996 41410
rect 8944 41346 8996 41352
rect 7564 41336 7616 41342
rect 7564 41278 7616 41284
rect 11716 41138 11744 480558
rect 14464 437504 14516 437510
rect 14464 437446 14516 437452
rect 13084 423700 13136 423706
rect 13084 423642 13136 423648
rect 12346 194576 12402 194585
rect 12346 194511 12402 194520
rect 12360 194426 12388 194511
rect 12530 194440 12586 194449
rect 12360 194398 12530 194426
rect 12530 194375 12586 194384
rect 13096 165578 13124 423642
rect 13084 165572 13136 165578
rect 13084 165514 13136 165520
rect 11704 41132 11756 41138
rect 11704 41074 11756 41080
rect 14476 39982 14504 437446
rect 14568 216646 14596 609962
rect 15844 552084 15896 552090
rect 15844 552026 15896 552032
rect 14556 216640 14608 216646
rect 14556 216582 14608 216588
rect 15856 168366 15884 552026
rect 24124 379568 24176 379574
rect 24124 379510 24176 379516
rect 22744 307828 22796 307834
rect 22744 307770 22796 307776
rect 22756 269822 22784 307770
rect 22744 269816 22796 269822
rect 22744 269758 22796 269764
rect 19984 267980 20036 267986
rect 19984 267922 20036 267928
rect 17224 266620 17276 266626
rect 17224 266562 17276 266568
rect 17236 237386 17264 266562
rect 17224 237380 17276 237386
rect 17224 237322 17276 237328
rect 19996 223514 20024 267922
rect 19984 223508 20036 223514
rect 19984 223450 20036 223456
rect 24136 200122 24164 379510
rect 24124 200116 24176 200122
rect 24124 200058 24176 200064
rect 22190 194576 22246 194585
rect 22190 194511 22246 194520
rect 27618 194576 27674 194585
rect 27618 194511 27620 194520
rect 22006 194440 22062 194449
rect 22204 194426 22232 194511
rect 27672 194511 27674 194520
rect 37188 194540 37240 194546
rect 27620 194482 27672 194488
rect 37188 194482 37240 194488
rect 22062 194398 22232 194426
rect 22006 194375 22062 194384
rect 37200 194313 37228 194482
rect 37186 194304 37242 194313
rect 37186 194239 37242 194248
rect 15844 168360 15896 168366
rect 15844 168302 15896 168308
rect 41340 42294 41368 700402
rect 89180 699718 89208 703520
rect 105464 700670 105492 703520
rect 111708 700732 111760 700738
rect 111708 700674 111760 700680
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 104808 700324 104860 700330
rect 104808 700266 104860 700272
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 60648 673532 60700 673538
rect 60648 673474 60700 673480
rect 51724 667956 51776 667962
rect 51724 667898 51776 667904
rect 41328 42288 41380 42294
rect 41328 42230 41380 42236
rect 51736 41954 51764 667898
rect 60556 368552 60608 368558
rect 60556 368494 60608 368500
rect 60464 272536 60516 272542
rect 60464 272478 60516 272484
rect 55864 268252 55916 268258
rect 55864 268194 55916 268200
rect 55128 266484 55180 266490
rect 55128 266426 55180 266432
rect 53748 266416 53800 266422
rect 53748 266358 53800 266364
rect 53656 263628 53708 263634
rect 53656 263570 53708 263576
rect 53564 220856 53616 220862
rect 53564 220798 53616 220804
rect 53472 216708 53524 216714
rect 53472 216650 53524 216656
rect 53380 205692 53432 205698
rect 53380 205634 53432 205640
rect 53288 193248 53340 193254
rect 53288 193190 53340 193196
rect 53196 180872 53248 180878
rect 53196 180814 53248 180820
rect 53104 135312 53156 135318
rect 53104 135254 53156 135260
rect 53116 42566 53144 135254
rect 53104 42560 53156 42566
rect 53104 42502 53156 42508
rect 51724 41948 51776 41954
rect 51724 41890 51776 41896
rect 14464 39976 14516 39982
rect 14464 39918 14516 39924
rect 53208 9178 53236 180814
rect 53196 9172 53248 9178
rect 53196 9114 53248 9120
rect 53300 9042 53328 193190
rect 53392 9314 53420 205634
rect 53380 9308 53432 9314
rect 53380 9250 53432 9256
rect 53288 9036 53340 9042
rect 53288 8978 53340 8984
rect 53484 8945 53512 216650
rect 53470 8936 53526 8945
rect 53470 8871 53526 8880
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 2976 7177 3004 7346
rect 2962 7168 3018 7177
rect 2962 7103 3018 7112
rect 53576 3738 53604 220798
rect 53668 6662 53696 263570
rect 53656 6656 53708 6662
rect 53656 6598 53708 6604
rect 53760 6458 53788 266358
rect 55036 263696 55088 263702
rect 55036 263638 55088 263644
rect 54944 213988 54996 213994
rect 54944 213930 54996 213936
rect 54852 202904 54904 202910
rect 54852 202846 54904 202852
rect 54760 128376 54812 128382
rect 54760 128318 54812 128324
rect 54668 120148 54720 120154
rect 54668 120090 54720 120096
rect 54680 9110 54708 120090
rect 54668 9104 54720 9110
rect 54772 9081 54800 128318
rect 54668 9046 54720 9052
rect 54758 9072 54814 9081
rect 54758 9007 54814 9016
rect 54864 6594 54892 202846
rect 54852 6588 54904 6594
rect 54852 6530 54904 6536
rect 53748 6452 53800 6458
rect 53748 6394 53800 6400
rect 54956 6254 54984 213930
rect 54944 6248 54996 6254
rect 54944 6190 54996 6196
rect 55048 4146 55076 263638
rect 55036 4140 55088 4146
rect 55036 4082 55088 4088
rect 53564 3732 53616 3738
rect 53564 3674 53616 3680
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 584 480 612 3470
rect 1688 480 1716 3470
rect 55140 3466 55168 266426
rect 55772 107704 55824 107710
rect 55772 107646 55824 107652
rect 55680 65340 55732 65346
rect 55680 65282 55732 65288
rect 55692 6526 55720 65282
rect 55784 42634 55812 107646
rect 55876 80034 55904 268194
rect 57704 267028 57756 267034
rect 57704 266970 57756 266976
rect 56324 266824 56376 266830
rect 56324 266766 56376 266772
rect 56232 266756 56284 266762
rect 56232 266698 56284 266704
rect 56140 212560 56192 212566
rect 56140 212502 56192 212508
rect 56048 117360 56100 117366
rect 56048 117302 56100 117308
rect 55956 100768 56008 100774
rect 55956 100710 56008 100716
rect 55864 80028 55916 80034
rect 55864 79970 55916 79976
rect 55864 74588 55916 74594
rect 55864 74530 55916 74536
rect 55772 42628 55824 42634
rect 55772 42570 55824 42576
rect 55876 6769 55904 74530
rect 55968 17950 55996 100710
rect 55956 17944 56008 17950
rect 55956 17886 56008 17892
rect 55862 6760 55918 6769
rect 55862 6695 55918 6704
rect 55680 6520 55732 6526
rect 55680 6462 55732 6468
rect 56060 6361 56088 117302
rect 56046 6352 56102 6361
rect 56046 6287 56102 6296
rect 56152 4049 56180 212502
rect 56244 42226 56272 266698
rect 56232 42220 56284 42226
rect 56232 42162 56284 42168
rect 56336 42158 56364 266766
rect 56508 263832 56560 263838
rect 56508 263774 56560 263780
rect 56416 263764 56468 263770
rect 56416 263706 56468 263712
rect 56324 42152 56376 42158
rect 56324 42094 56376 42100
rect 56138 4040 56194 4049
rect 56428 4010 56456 263706
rect 56138 3975 56194 3984
rect 56416 4004 56468 4010
rect 56416 3946 56468 3952
rect 55128 3460 55180 3466
rect 55128 3402 55180 3408
rect 56520 3330 56548 263774
rect 57612 182232 57664 182238
rect 57612 182174 57664 182180
rect 57520 175296 57572 175302
rect 57520 175238 57572 175244
rect 57428 142656 57480 142662
rect 57428 142598 57480 142604
rect 57334 142080 57390 142089
rect 57334 142015 57390 142024
rect 57244 129804 57296 129810
rect 57244 129746 57296 129752
rect 57152 111852 57204 111858
rect 57152 111794 57204 111800
rect 57060 43444 57112 43450
rect 57060 43386 57112 43392
rect 57072 41206 57100 43386
rect 57060 41200 57112 41206
rect 57060 41142 57112 41148
rect 57164 3874 57192 111794
rect 57256 6225 57284 129746
rect 57242 6216 57298 6225
rect 57242 6151 57298 6160
rect 57152 3868 57204 3874
rect 57152 3810 57204 3816
rect 57348 3505 57376 142015
rect 57334 3496 57390 3505
rect 57334 3431 57390 3440
rect 57440 3369 57468 142598
rect 57532 17406 57560 175238
rect 57520 17400 57572 17406
rect 57520 17342 57572 17348
rect 57624 3806 57652 182174
rect 57612 3800 57664 3806
rect 57612 3742 57664 3748
rect 57716 3670 57744 266970
rect 57796 266960 57848 266966
rect 57796 266902 57848 266908
rect 57808 4078 57836 266902
rect 57888 266892 57940 266898
rect 57888 266834 57940 266840
rect 57796 4072 57848 4078
rect 57796 4014 57848 4020
rect 57900 3942 57928 266834
rect 60280 262812 60332 262818
rect 60280 262754 60332 262760
rect 59360 260840 59412 260846
rect 59360 260782 59412 260788
rect 59372 260409 59400 260782
rect 59358 260400 59414 260409
rect 59358 260335 59414 260344
rect 59266 240000 59322 240009
rect 59266 239935 59322 239944
rect 59174 234016 59230 234025
rect 59174 233951 59230 233960
rect 59082 229664 59138 229673
rect 59082 229599 59138 229608
rect 58898 187232 58954 187241
rect 58898 187167 58954 187176
rect 58806 174176 58862 174185
rect 58806 174111 58862 174120
rect 58714 146432 58770 146441
rect 58714 146367 58770 146376
rect 58532 131164 58584 131170
rect 58532 131106 58584 131112
rect 58440 122936 58492 122942
rect 58440 122878 58492 122884
rect 58452 36650 58480 122878
rect 58440 36644 58492 36650
rect 58440 36586 58492 36592
rect 58544 31210 58572 131106
rect 58622 120048 58678 120057
rect 58622 119983 58678 119992
rect 58532 31204 58584 31210
rect 58532 31146 58584 31152
rect 58636 11762 58664 119983
rect 58728 26994 58756 146367
rect 58820 35358 58848 174111
rect 58808 35352 58860 35358
rect 58808 35294 58860 35300
rect 58912 35290 58940 187167
rect 58990 185872 59046 185881
rect 58990 185807 59046 185816
rect 58900 35284 58952 35290
rect 58900 35226 58952 35232
rect 58716 26988 58768 26994
rect 58716 26930 58768 26936
rect 59004 18630 59032 185807
rect 59096 31074 59124 229599
rect 59084 31068 59136 31074
rect 59084 31010 59136 31016
rect 59188 24206 59216 233951
rect 59176 24200 59228 24206
rect 59176 24142 59228 24148
rect 58992 18624 59044 18630
rect 58992 18566 59044 18572
rect 59280 16046 59308 239935
rect 59360 223576 59412 223582
rect 59360 223518 59412 223524
rect 59372 222329 59400 223518
rect 59358 222320 59414 222329
rect 59358 222255 59414 222264
rect 59358 220960 59414 220969
rect 59358 220895 59414 220904
rect 59372 220862 59400 220895
rect 59360 220856 59412 220862
rect 59360 220798 59412 220804
rect 59450 217968 59506 217977
rect 59450 217903 59506 217912
rect 59464 216714 59492 217903
rect 59452 216708 59504 216714
rect 59452 216650 59504 216656
rect 59360 216640 59412 216646
rect 59358 216608 59360 216617
rect 59412 216608 59414 216617
rect 59358 216543 59414 216552
rect 59358 214976 59414 214985
rect 59358 214911 59414 214920
rect 59372 213994 59400 214911
rect 59360 213988 59412 213994
rect 59360 213930 59412 213936
rect 59358 213616 59414 213625
rect 59358 213551 59414 213560
rect 59372 212566 59400 213551
rect 59360 212560 59412 212566
rect 59360 212502 59412 212508
rect 59358 206272 59414 206281
rect 59358 206207 59414 206216
rect 59372 205698 59400 206207
rect 59360 205692 59412 205698
rect 59360 205634 59412 205640
rect 59358 203280 59414 203289
rect 59358 203215 59414 203224
rect 59372 202910 59400 203215
rect 59360 202904 59412 202910
rect 59360 202846 59412 202852
rect 59360 200116 59412 200122
rect 59360 200058 59412 200064
rect 59372 198937 59400 200058
rect 59358 198928 59414 198937
rect 59358 198863 59414 198872
rect 59358 194576 59414 194585
rect 59358 194511 59414 194520
rect 59372 193254 59400 194511
rect 59360 193248 59412 193254
rect 59360 193190 59412 193196
rect 60292 190233 60320 262754
rect 60476 257417 60504 272478
rect 60462 257408 60518 257417
rect 60462 257343 60518 257352
rect 60462 237008 60518 237017
rect 60462 236943 60518 236952
rect 60370 193216 60426 193225
rect 60370 193151 60426 193160
rect 60278 190224 60334 190233
rect 60278 190159 60334 190168
rect 59360 189032 59412 189038
rect 59360 188974 59412 188980
rect 59372 188873 59400 188974
rect 59358 188864 59414 188873
rect 59358 188799 59414 188808
rect 59910 182880 59966 182889
rect 59910 182815 59966 182824
rect 59924 182238 59952 182815
rect 59912 182232 59964 182238
rect 59912 182174 59964 182180
rect 59358 181520 59414 181529
rect 59358 181455 59414 181464
rect 59372 180878 59400 181455
rect 59360 180872 59412 180878
rect 59360 180814 59412 180820
rect 59542 175536 59598 175545
rect 59542 175471 59598 175480
rect 59556 175302 59584 175471
rect 59544 175296 59596 175302
rect 59544 175238 59596 175244
rect 59360 168360 59412 168366
rect 59360 168302 59412 168308
rect 59372 168201 59400 168302
rect 59358 168192 59414 168201
rect 59358 168127 59414 168136
rect 59360 165572 59412 165578
rect 59360 165514 59412 165520
rect 59372 165481 59400 165514
rect 59358 165472 59414 165481
rect 59358 165407 59414 165416
rect 60094 153776 60150 153785
rect 60094 153711 60150 153720
rect 59358 150784 59414 150793
rect 59358 150719 59414 150728
rect 59372 150482 59400 150719
rect 59360 150476 59412 150482
rect 59360 150418 59412 150424
rect 59358 143440 59414 143449
rect 59358 143375 59414 143384
rect 59372 142662 59400 143375
rect 59360 142656 59412 142662
rect 59360 142598 59412 142604
rect 59358 131744 59414 131753
rect 59358 131679 59414 131688
rect 59372 131170 59400 131679
rect 59360 131164 59412 131170
rect 59360 131106 59412 131112
rect 59726 130384 59782 130393
rect 59726 130319 59782 130328
rect 59740 129810 59768 130319
rect 59728 129804 59780 129810
rect 59728 129746 59780 129752
rect 59358 128752 59414 128761
rect 59358 128687 59414 128696
rect 59372 128382 59400 128687
rect 59360 128376 59412 128382
rect 59360 128318 59412 128324
rect 59358 121408 59414 121417
rect 59358 121343 59414 121352
rect 59372 120154 59400 121343
rect 59360 120148 59412 120154
rect 59360 120090 59412 120096
rect 59358 118688 59414 118697
rect 59358 118623 59414 118632
rect 59372 117366 59400 118623
rect 59360 117360 59412 117366
rect 59360 117302 59412 117308
rect 59634 112704 59690 112713
rect 59634 112639 59690 112648
rect 59648 111858 59676 112639
rect 59636 111852 59688 111858
rect 59636 111794 59688 111800
rect 59358 104000 59414 104009
rect 59358 103935 59414 103944
rect 59372 103562 59400 103935
rect 59360 103556 59412 103562
rect 59360 103498 59412 103504
rect 59358 101008 59414 101017
rect 59358 100943 59414 100952
rect 59372 100774 59400 100943
rect 59360 100768 59412 100774
rect 59360 100710 59412 100716
rect 60108 98938 60136 153711
rect 60186 133104 60242 133113
rect 60186 133039 60242 133048
rect 60096 98932 60148 98938
rect 60096 98874 60148 98880
rect 59360 91044 59412 91050
rect 59360 90986 59412 90992
rect 59372 90953 59400 90986
rect 59358 90944 59414 90953
rect 59358 90879 59414 90888
rect 59726 87952 59782 87961
rect 59726 87887 59782 87896
rect 59634 83600 59690 83609
rect 59634 83535 59690 83544
rect 59360 78668 59412 78674
rect 59360 78610 59412 78616
rect 59372 77625 59400 78610
rect 59358 77616 59414 77625
rect 59358 77551 59414 77560
rect 59358 74624 59414 74633
rect 59358 74559 59360 74568
rect 59412 74559 59414 74568
rect 59360 74530 59412 74536
rect 59358 65920 59414 65929
rect 59358 65855 59414 65864
rect 59372 65346 59400 65855
rect 59360 65340 59412 65346
rect 59360 65282 59412 65288
rect 59360 60716 59412 60722
rect 59360 60658 59412 60664
rect 59372 60217 59400 60658
rect 59358 60208 59414 60217
rect 59358 60143 59414 60152
rect 59648 37942 59676 83535
rect 59740 39370 59768 87887
rect 60200 81569 60228 133039
rect 60278 123040 60334 123049
rect 60278 122975 60334 122984
rect 60292 122942 60320 122975
rect 60280 122936 60332 122942
rect 60280 122878 60332 122884
rect 60278 105360 60334 105369
rect 60278 105295 60334 105304
rect 60186 81560 60242 81569
rect 60186 81495 60242 81504
rect 60002 80608 60058 80617
rect 60002 80543 60058 80552
rect 59910 64560 59966 64569
rect 59910 64495 59966 64504
rect 59728 39364 59780 39370
rect 59728 39306 59780 39312
rect 59636 37936 59688 37942
rect 59636 37878 59688 37884
rect 59924 33862 59952 64495
rect 60016 43586 60044 80543
rect 60094 79248 60150 79257
rect 60094 79183 60150 79192
rect 60004 43580 60056 43586
rect 60004 43522 60056 43528
rect 60108 36582 60136 79183
rect 60292 43518 60320 105295
rect 60280 43512 60332 43518
rect 60280 43454 60332 43460
rect 60384 42974 60412 193151
rect 60476 75857 60504 236943
rect 60568 149433 60596 368494
rect 60660 172825 60688 673474
rect 73068 592068 73120 592074
rect 73068 592010 73120 592016
rect 62488 438932 62540 438938
rect 62488 438874 62540 438880
rect 61200 310548 61252 310554
rect 61200 310490 61252 310496
rect 60924 271176 60976 271182
rect 60924 271118 60976 271124
rect 60738 253056 60794 253065
rect 60738 252991 60794 253000
rect 60646 172816 60702 172825
rect 60646 172751 60702 172760
rect 60554 149424 60610 149433
rect 60554 149359 60610 149368
rect 60648 128376 60700 128382
rect 60648 128318 60700 128324
rect 60660 111353 60688 128318
rect 60646 111344 60702 111353
rect 60646 111279 60702 111288
rect 60646 106992 60702 107001
rect 60646 106927 60702 106936
rect 60554 97744 60610 97753
rect 60554 97679 60610 97688
rect 60462 75848 60518 75857
rect 60462 75783 60518 75792
rect 60462 49600 60518 49609
rect 60462 49535 60518 49544
rect 60476 43858 60504 49535
rect 60464 43852 60516 43858
rect 60464 43794 60516 43800
rect 60372 42968 60424 42974
rect 60372 42910 60424 42916
rect 60096 36576 60148 36582
rect 60096 36518 60148 36524
rect 59912 33856 59964 33862
rect 59912 33798 59964 33804
rect 60568 28422 60596 97679
rect 60556 28416 60608 28422
rect 60556 28358 60608 28364
rect 59268 16040 59320 16046
rect 59268 15982 59320 15988
rect 58624 11756 58676 11762
rect 58624 11698 58676 11704
rect 60660 10334 60688 106927
rect 60752 11830 60780 252991
rect 60830 250064 60886 250073
rect 60830 249999 60886 250008
rect 60844 22846 60872 249999
rect 60936 238377 60964 271118
rect 61014 251696 61070 251705
rect 61014 251631 61070 251640
rect 60922 238368 60978 238377
rect 60922 238303 60978 238312
rect 60922 219600 60978 219609
rect 60922 219535 60978 219544
rect 60936 39438 60964 219535
rect 61028 73137 61056 251631
rect 61106 248704 61162 248713
rect 61106 248639 61162 248648
rect 61120 208321 61148 248639
rect 61106 208312 61162 208321
rect 61106 208247 61162 208256
rect 61106 163840 61162 163849
rect 61106 163775 61162 163784
rect 61014 73128 61070 73137
rect 61014 73063 61070 73072
rect 61014 70272 61070 70281
rect 61014 70207 61070 70216
rect 61028 43790 61056 70207
rect 61016 43784 61068 43790
rect 61016 43726 61068 43732
rect 60924 39432 60976 39438
rect 60924 39374 60976 39380
rect 60832 22840 60884 22846
rect 60832 22782 60884 22788
rect 60740 11824 60792 11830
rect 60740 11766 60792 11772
rect 60648 10328 60700 10334
rect 60648 10270 60700 10276
rect 61120 7818 61148 163775
rect 61212 159497 61240 310490
rect 61290 223952 61346 223961
rect 61290 223887 61346 223896
rect 61304 193361 61332 223887
rect 62394 205864 62450 205873
rect 62394 205799 62450 205808
rect 62408 201521 62436 205799
rect 62394 201512 62450 201521
rect 62394 201447 62450 201456
rect 61290 193352 61346 193361
rect 61290 193287 61346 193296
rect 61290 191584 61346 191593
rect 61290 191519 61346 191528
rect 61198 159488 61254 159497
rect 61198 159423 61254 159432
rect 61198 94752 61254 94761
rect 61198 94687 61254 94696
rect 61212 25634 61240 94687
rect 61304 43722 61332 191519
rect 62396 128376 62448 128382
rect 62500 128364 62528 438874
rect 64052 270632 64104 270638
rect 64052 270574 64104 270580
rect 64064 264996 64092 270574
rect 69020 268184 69072 268190
rect 69020 268126 69072 268132
rect 67916 266688 67968 266694
rect 67916 266630 67968 266636
rect 66996 266484 67048 266490
rect 66996 266426 67048 266432
rect 65892 266416 65944 266422
rect 65892 266358 65944 266364
rect 64970 265432 65026 265441
rect 64970 265367 65026 265376
rect 64984 264996 65012 265367
rect 65904 264996 65932 266358
rect 67008 264996 67036 266426
rect 67928 264996 67956 266630
rect 69032 266354 69060 268126
rect 71964 266484 72016 266490
rect 71964 266426 72016 266432
rect 69020 266348 69072 266354
rect 69020 266290 69072 266296
rect 68836 265124 68888 265130
rect 68836 265066 68888 265072
rect 68848 264996 68876 265066
rect 71976 264996 72004 266426
rect 73080 265010 73108 592010
rect 89640 278050 89668 699654
rect 100668 451308 100720 451314
rect 100668 451250 100720 451256
rect 89628 278044 89680 278050
rect 89628 277986 89680 277992
rect 98644 270700 98696 270706
rect 98644 270642 98696 270648
rect 73804 270564 73856 270570
rect 73804 270506 73856 270512
rect 72910 264982 73108 265010
rect 73816 264996 73844 270506
rect 97540 270020 97592 270026
rect 97540 269962 97592 269968
rect 76748 269816 76800 269822
rect 76748 269758 76800 269764
rect 74906 269240 74962 269249
rect 74906 269175 74962 269184
rect 74920 264996 74948 269175
rect 76760 264996 76788 269758
rect 86682 268424 86738 268433
rect 86682 268359 86738 268368
rect 78770 267200 78826 267209
rect 78770 267135 78826 267144
rect 78784 264996 78812 267135
rect 84660 267096 84712 267102
rect 84660 267038 84712 267044
rect 79874 265296 79930 265305
rect 79874 265231 79930 265240
rect 79888 264996 79916 265231
rect 84672 264996 84700 267038
rect 86696 264996 86724 268359
rect 89628 267368 89680 267374
rect 89628 267310 89680 267316
rect 88706 265840 88762 265849
rect 88706 265775 88762 265784
rect 88720 264996 88748 265775
rect 89640 264996 89668 267310
rect 96620 265328 96672 265334
rect 96620 265270 96672 265276
rect 96632 264996 96660 265270
rect 97552 264996 97580 269962
rect 98656 264996 98684 270642
rect 100680 267714 100708 451250
rect 102506 267880 102562 267889
rect 102506 267815 102562 267824
rect 99564 267708 99616 267714
rect 99564 267650 99616 267656
rect 100668 267708 100720 267714
rect 100668 267650 100720 267656
rect 99576 264996 99604 267650
rect 102520 264996 102548 267815
rect 103610 266792 103666 266801
rect 103610 266727 103666 266736
rect 103624 264996 103652 266727
rect 104820 265010 104848 700266
rect 111720 267714 111748 700674
rect 137848 700602 137876 703520
rect 154132 700738 154160 703520
rect 154120 700732 154172 700738
rect 154120 700674 154172 700680
rect 169760 700664 169812 700670
rect 169760 700606 169812 700612
rect 137836 700596 137888 700602
rect 137836 700538 137888 700544
rect 143448 700460 143500 700466
rect 143448 700402 143500 700408
rect 120356 269952 120408 269958
rect 120356 269894 120408 269900
rect 112444 269272 112496 269278
rect 112444 269214 112496 269220
rect 110420 267708 110472 267714
rect 110420 267650 110472 267656
rect 111708 267708 111760 267714
rect 111708 267650 111760 267656
rect 107474 266928 107530 266937
rect 107474 266863 107530 266872
rect 106554 266520 106610 266529
rect 106554 266455 106610 266464
rect 104558 264982 104848 265010
rect 106568 264996 106596 266455
rect 107488 264996 107516 266863
rect 110432 264996 110460 267650
rect 112456 264996 112484 269214
rect 115388 267232 115440 267238
rect 115388 267174 115440 267180
rect 114466 265160 114522 265169
rect 114466 265095 114522 265104
rect 114480 264996 114508 265095
rect 115400 264996 115428 267174
rect 116308 267028 116360 267034
rect 116308 266970 116360 266976
rect 116320 264996 116348 266970
rect 117412 266620 117464 266626
rect 117412 266562 117464 266568
rect 117424 264996 117452 266562
rect 120368 264996 120396 269894
rect 139124 269408 139176 269414
rect 139124 269350 139176 269356
rect 128268 266960 128320 266966
rect 128268 266902 128320 266908
rect 132868 266960 132920 266966
rect 132868 266902 132920 266908
rect 126980 266688 127032 266694
rect 126980 266630 127032 266636
rect 124220 266620 124272 266626
rect 124220 266562 124272 266568
rect 122380 266416 122432 266422
rect 122380 266358 122432 266364
rect 122392 264996 122420 266358
rect 124232 264996 124260 266562
rect 126992 265577 127020 266630
rect 126978 265568 127034 265577
rect 126978 265503 127034 265512
rect 128280 264996 128308 266902
rect 129186 266520 129242 266529
rect 129186 266455 129242 266464
rect 128360 266416 128412 266422
rect 128360 266358 128412 266364
rect 128372 265674 128400 266358
rect 128360 265668 128412 265674
rect 128360 265610 128412 265616
rect 129200 264996 129228 266455
rect 132880 264450 132908 266902
rect 137100 266892 137152 266898
rect 137100 266834 137152 266840
rect 137112 264996 137140 266834
rect 139136 264996 139164 269350
rect 142066 266656 142122 266665
rect 142066 266591 142122 266600
rect 142080 264996 142108 266591
rect 143460 265010 143488 700402
rect 160008 462392 160060 462398
rect 160008 462334 160060 462340
rect 156972 269680 157024 269686
rect 156972 269622 157024 269628
rect 152924 269612 152976 269618
rect 152924 269554 152976 269560
rect 145012 267844 145064 267850
rect 145012 267786 145064 267792
rect 143198 264982 143488 265010
rect 145024 264996 145052 267786
rect 149058 266928 149114 266937
rect 149058 266863 149114 266872
rect 149072 264996 149100 266863
rect 149980 265396 150032 265402
rect 149980 265338 150032 265344
rect 149992 264996 150020 265338
rect 152936 264996 152964 269554
rect 154948 266824 155000 266830
rect 154948 266766 155000 266772
rect 154960 264996 154988 266766
rect 155868 265872 155920 265878
rect 155868 265814 155920 265820
rect 155880 264996 155908 265814
rect 156984 264996 157012 269622
rect 157892 266552 157944 266558
rect 157892 266494 157944 266500
rect 157904 264996 157932 266494
rect 160020 266422 160048 462334
rect 164884 269748 164936 269754
rect 164884 269690 164936 269696
rect 163964 269340 164016 269346
rect 163964 269282 164016 269288
rect 163044 268660 163096 268666
rect 163044 268602 163096 268608
rect 158996 266416 159048 266422
rect 158996 266358 159048 266364
rect 160008 266416 160060 266422
rect 160008 266358 160060 266364
rect 159008 264996 159036 266358
rect 161940 265192 161992 265198
rect 161940 265134 161992 265140
rect 161952 264996 161980 265134
rect 163056 265010 163084 268602
rect 163412 266416 163464 266422
rect 163412 266358 163464 266364
rect 162886 264982 163084 265010
rect 161112 264512 161164 264518
rect 160862 264460 161112 264466
rect 160862 264454 161164 264460
rect 132868 264444 132920 264450
rect 160862 264438 161152 264454
rect 132868 264386 132920 264392
rect 136456 264376 136508 264382
rect 63222 264344 63278 264353
rect 62974 264302 63222 264330
rect 113546 264344 113602 264353
rect 81452 264314 81742 264330
rect 85592 264314 85790 264330
rect 87432 264314 87814 264330
rect 63222 264279 63278 264288
rect 81440 264308 81742 264314
rect 81492 264302 81742 264308
rect 85580 264308 85790 264314
rect 81440 264250 81492 264256
rect 85632 264302 85790 264308
rect 87420 264308 87814 264314
rect 85580 264250 85632 264256
rect 87472 264302 87814 264308
rect 108422 264314 108712 264330
rect 108422 264308 108724 264314
rect 108422 264302 108672 264308
rect 87420 264250 87472 264256
rect 113390 264302 113546 264330
rect 132158 264314 132356 264330
rect 133262 264314 133552 264330
rect 134182 264314 134472 264330
rect 136206 264324 136456 264330
rect 163424 264353 163452 266358
rect 163976 264996 164004 269282
rect 164148 266824 164200 266830
rect 164148 266766 164200 266772
rect 164160 265742 164188 266766
rect 164148 265736 164200 265742
rect 164148 265678 164200 265684
rect 164896 264996 164924 269690
rect 168748 268048 168800 268054
rect 168748 267990 168800 267996
rect 168760 264996 168788 267990
rect 169772 265146 169800 700606
rect 170324 700505 170352 703520
rect 170310 700496 170366 700505
rect 170310 700431 170366 700440
rect 190460 594856 190512 594862
rect 190460 594798 190512 594804
rect 183560 365764 183612 365770
rect 183560 365706 183612 365712
rect 181628 269544 181680 269550
rect 181628 269486 181680 269492
rect 174820 269476 174872 269482
rect 174820 269418 174872 269424
rect 172796 268456 172848 268462
rect 172796 268398 172848 268404
rect 171876 265260 171928 265266
rect 171876 265202 171928 265208
rect 169772 265118 170444 265146
rect 170416 265010 170444 265118
rect 170416 264982 170798 265010
rect 171888 264996 171916 265202
rect 172808 264996 172836 268398
rect 174832 264996 174860 269418
rect 178684 268388 178736 268394
rect 178684 268330 178736 268336
rect 178696 264996 178724 268330
rect 180708 266960 180760 266966
rect 180708 266902 180760 266908
rect 179788 266756 179840 266762
rect 179788 266698 179840 266704
rect 179800 264996 179828 266698
rect 180720 264996 180748 266902
rect 181640 264996 181668 269486
rect 183572 265010 183600 365706
rect 189540 269884 189592 269890
rect 189540 269826 189592 269832
rect 187700 269816 187752 269822
rect 187700 269758 187752 269764
rect 183572 264982 183678 265010
rect 187712 264996 187740 269758
rect 188620 267912 188672 267918
rect 188620 267854 188672 267860
rect 188632 264996 188660 267854
rect 189552 264996 189580 269826
rect 190472 265146 190500 594798
rect 202800 273970 202828 703520
rect 218992 700369 219020 703520
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 235908 700664 235960 700670
rect 235908 700606 235960 700612
rect 218978 700360 219034 700369
rect 218978 700295 219034 700304
rect 223488 603152 223540 603158
rect 223488 603094 223540 603100
rect 205640 495508 205692 495514
rect 205640 495450 205692 495456
rect 202788 273964 202840 273970
rect 202788 273906 202840 273912
rect 199474 269376 199530 269385
rect 199474 269311 199530 269320
rect 197452 266824 197504 266830
rect 197452 266766 197504 266772
rect 198556 266824 198608 266830
rect 198556 266766 198608 266772
rect 194508 266756 194560 266762
rect 194508 266698 194560 266704
rect 190472 265118 190960 265146
rect 190932 264874 190960 265118
rect 194520 264996 194548 266698
rect 197464 264996 197492 266766
rect 198568 264996 198596 266766
rect 199488 264996 199516 269311
rect 200394 268016 200450 268025
rect 200394 267951 200450 267960
rect 200408 264996 200436 267951
rect 205652 267458 205680 495450
rect 216588 298172 216640 298178
rect 216588 298114 216640 298120
rect 211436 268524 211488 268530
rect 211436 268466 211488 268472
rect 205652 267430 206140 267458
rect 206112 265010 206140 267430
rect 210332 266416 210384 266422
rect 210332 266358 210384 266364
rect 206112 264982 206494 265010
rect 210344 264996 210372 266358
rect 211448 264996 211476 268466
rect 213276 268320 213328 268326
rect 213276 268262 213328 268268
rect 213288 264996 213316 268262
rect 214380 268252 214432 268258
rect 214380 268194 214432 268200
rect 214392 264996 214420 268194
rect 215300 265532 215352 265538
rect 215300 265474 215352 265480
rect 215312 264996 215340 265474
rect 216600 265010 216628 298114
rect 220268 268592 220320 268598
rect 220268 268534 220320 268540
rect 216246 264982 216628 265010
rect 220280 264996 220308 268534
rect 221188 265464 221240 265470
rect 221188 265406 221240 265412
rect 221200 264996 221228 265406
rect 223500 265010 223528 603094
rect 235920 461650 235948 700606
rect 253940 700392 253992 700398
rect 267660 700369 267688 703520
rect 283012 700596 283064 700602
rect 283012 700538 283064 700544
rect 269120 700528 269172 700534
rect 269120 700470 269172 700476
rect 253940 700334 253992 700340
rect 267646 700360 267702 700369
rect 249708 532772 249760 532778
rect 249708 532714 249760 532720
rect 242900 509312 242952 509318
rect 242900 509254 242952 509260
rect 235908 461644 235960 461650
rect 235908 461586 235960 461592
rect 242912 268818 242940 509254
rect 246026 269648 246082 269657
rect 246026 269583 246082 269592
rect 244922 269512 244978 269521
rect 244922 269447 244978 269456
rect 242912 268790 243676 268818
rect 236092 268252 236144 268258
rect 236092 268194 236144 268200
rect 229100 267980 229152 267986
rect 229100 267922 229152 267928
rect 230204 267980 230256 267986
rect 230204 267922 230256 267928
rect 226156 266892 226208 266898
rect 226156 266834 226208 266840
rect 223238 264982 223528 265010
rect 226168 264996 226196 266834
rect 226248 266416 226300 266422
rect 226248 266358 226300 266364
rect 190932 264846 191590 264874
rect 209686 264480 209742 264489
rect 208334 264450 208440 264466
rect 208334 264444 208452 264450
rect 208334 264438 208400 264444
rect 209438 264438 209686 264466
rect 209686 264415 209742 264424
rect 208400 264386 208452 264392
rect 226260 264382 226288 266358
rect 229112 264996 229140 267922
rect 230216 264996 230244 267922
rect 231124 265804 231176 265810
rect 231124 265746 231176 265752
rect 231136 264996 231164 265746
rect 233056 265056 233108 265062
rect 233108 265004 233174 265010
rect 233056 264998 233174 265004
rect 233068 264982 233174 264998
rect 236104 264996 236132 268194
rect 238114 267064 238170 267073
rect 238114 266999 238170 267008
rect 237012 266960 237064 266966
rect 237012 266902 237064 266908
rect 237024 264996 237052 266902
rect 238128 264996 238156 266999
rect 241058 265704 241114 265713
rect 241058 265639 241114 265648
rect 241072 264996 241100 265639
rect 243648 265010 243676 268790
rect 243648 264982 244030 265010
rect 244936 264996 244964 269447
rect 246040 264996 246068 269583
rect 249720 267714 249748 532714
rect 252836 267776 252888 267782
rect 252836 267718 252888 267724
rect 248972 267708 249024 267714
rect 248972 267650 249024 267656
rect 249708 267708 249760 267714
rect 249708 267650 249760 267656
rect 248984 264996 249012 267650
rect 249892 267164 249944 267170
rect 249892 267106 249944 267112
rect 249904 264996 249932 267106
rect 252848 264996 252876 267718
rect 253952 264996 253980 700334
rect 267646 700295 267702 700304
rect 255320 567248 255372 567254
rect 255320 567190 255372 567196
rect 255332 265010 255360 567190
rect 262772 269204 262824 269210
rect 262772 269146 262824 269152
rect 260748 269136 260800 269142
rect 260748 269078 260800 269084
rect 259828 267300 259880 267306
rect 259828 267242 259880 267248
rect 257988 267232 258040 267238
rect 257988 267174 258040 267180
rect 256884 266688 256936 266694
rect 256884 266630 256936 266636
rect 255332 264982 255806 265010
rect 256896 264996 256924 266630
rect 257802 266384 257858 266393
rect 257802 266319 257858 266328
rect 257816 264996 257844 266319
rect 258000 265742 258028 267174
rect 259460 266484 259512 266490
rect 259460 266426 259512 266432
rect 257988 265736 258040 265742
rect 257988 265678 258040 265684
rect 251942 264586 252232 264602
rect 258934 264586 259224 264602
rect 251942 264580 252244 264586
rect 251942 264574 252192 264580
rect 258934 264580 259236 264586
rect 258934 264574 259184 264580
rect 252192 264522 252244 264528
rect 259184 264522 259236 264528
rect 226248 264376 226300 264382
rect 159546 264344 159602 264353
rect 136206 264318 136508 264324
rect 132158 264308 132368 264314
rect 132158 264302 132316 264308
rect 113546 264279 113602 264288
rect 108672 264250 108724 264256
rect 133262 264308 133564 264314
rect 133262 264302 133512 264308
rect 132316 264250 132368 264256
rect 134182 264308 134484 264314
rect 134182 264302 134432 264308
rect 133512 264250 133564 264256
rect 136206 264302 136496 264318
rect 144118 264314 144408 264330
rect 147692 264314 147982 264330
rect 144118 264308 144420 264314
rect 144118 264302 144368 264308
rect 134432 264250 134484 264256
rect 144368 264250 144420 264256
rect 147680 264308 147982 264314
rect 147732 264302 147982 264308
rect 163410 264344 163466 264353
rect 159602 264302 159942 264330
rect 159546 264279 159602 264288
rect 201682 264344 201738 264353
rect 173742 264314 173848 264330
rect 173742 264308 173860 264314
rect 173742 264302 173808 264308
rect 163410 264279 163466 264288
rect 147680 264250 147732 264256
rect 201526 264302 201682 264330
rect 222566 264344 222622 264353
rect 202446 264314 202736 264330
rect 218270 264314 218560 264330
rect 202446 264308 202748 264314
rect 202446 264302 202696 264308
rect 201682 264279 201738 264288
rect 173808 264250 173860 264256
rect 218270 264308 218572 264314
rect 218270 264302 218520 264308
rect 202696 264250 202748 264256
rect 222318 264302 222566 264330
rect 224158 264314 224448 264330
rect 242256 264376 242308 264382
rect 226248 264318 226300 264324
rect 242006 264324 242256 264330
rect 259472 264353 259500 266426
rect 259840 264996 259868 267242
rect 260760 264996 260788 269078
rect 262784 264996 262812 269146
rect 264794 267336 264850 267345
rect 264794 267271 264850 267280
rect 263692 267232 263744 267238
rect 263692 267174 263744 267180
rect 263598 266656 263654 266665
rect 263598 266591 263654 266600
rect 263612 266354 263640 266591
rect 263600 266348 263652 266354
rect 263600 266290 263652 266296
rect 263704 264996 263732 267174
rect 264808 264996 264836 267271
rect 265716 267028 265768 267034
rect 265716 266970 265768 266976
rect 265728 264996 265756 266970
rect 267740 266484 267792 266490
rect 267740 266426 267792 266432
rect 267752 264996 267780 266426
rect 268686 264994 268976 265010
rect 268686 264988 268988 264994
rect 268686 264982 268936 264988
rect 268936 264930 268988 264936
rect 269132 264874 269160 700470
rect 282920 692844 282972 692850
rect 282920 692786 282972 692792
rect 281448 545148 281500 545154
rect 281448 545090 281500 545096
rect 273628 268116 273680 268122
rect 273628 268058 273680 268064
rect 270500 267368 270552 267374
rect 270500 267310 270552 267316
rect 270512 266665 270540 267310
rect 270498 266656 270554 266665
rect 270498 266591 270554 266600
rect 270684 266552 270736 266558
rect 270684 266494 270736 266500
rect 270696 264996 270724 266494
rect 271786 266384 271842 266393
rect 271786 266319 271842 266328
rect 271800 266286 271828 266319
rect 271788 266280 271840 266286
rect 271788 266222 271840 266228
rect 271786 265024 271842 265033
rect 271630 264982 271786 265010
rect 273640 264996 273668 268058
rect 281460 267714 281488 545090
rect 281540 461644 281592 461650
rect 281540 461586 281592 461592
rect 280620 267708 280672 267714
rect 280620 267650 280672 267656
rect 281448 267708 281500 267714
rect 281448 267650 281500 267656
rect 277676 266416 277728 266422
rect 277676 266358 277728 266364
rect 275652 265600 275704 265606
rect 275652 265542 275704 265548
rect 275664 264996 275692 265542
rect 277688 264996 277716 266358
rect 280632 264996 280660 267650
rect 281356 267300 281408 267306
rect 281356 267242 281408 267248
rect 281078 267064 281134 267073
rect 281078 266999 281134 267008
rect 281172 267028 281224 267034
rect 280896 266416 280948 266422
rect 280896 266358 280948 266364
rect 271786 264959 271842 264968
rect 269132 264846 269790 264874
rect 268290 264616 268346 264625
rect 268290 264551 268346 264560
rect 279882 264616 279938 264625
rect 279882 264551 279938 264560
rect 268304 264353 268332 264551
rect 279896 264353 279924 264551
rect 255134 264344 255190 264353
rect 242006 264318 242308 264324
rect 224158 264308 224460 264314
rect 224158 264302 224408 264308
rect 222566 264279 222622 264288
rect 218520 264250 218572 264256
rect 242006 264302 242296 264318
rect 254886 264302 255134 264330
rect 255134 264279 255190 264288
rect 259458 264344 259514 264353
rect 259458 264279 259514 264288
rect 268290 264344 268346 264353
rect 275006 264344 275062 264353
rect 274758 264302 275006 264330
rect 268290 264279 268346 264288
rect 279882 264344 279938 264353
rect 278622 264314 278728 264330
rect 279542 264314 279832 264330
rect 278622 264308 278740 264314
rect 278622 264302 278688 264308
rect 275006 264279 275062 264288
rect 224408 264250 224460 264256
rect 279542 264308 279844 264314
rect 279542 264302 279792 264308
rect 278688 264250 278740 264256
rect 279882 264279 279938 264288
rect 280804 264308 280856 264314
rect 279792 264250 279844 264256
rect 280804 264250 280856 264256
rect 280816 253230 280844 264250
rect 280908 260234 280936 266358
rect 280986 263528 281042 263537
rect 280986 263463 281042 263472
rect 281000 263226 281028 263463
rect 280988 263220 281040 263226
rect 280988 263162 281040 263168
rect 281092 263106 281120 266999
rect 281172 266970 281224 266976
rect 281000 263078 281120 263106
rect 281000 261526 281028 263078
rect 281080 263016 281132 263022
rect 281080 262958 281132 262964
rect 280988 261520 281040 261526
rect 280988 261462 281040 261468
rect 280896 260228 280948 260234
rect 280896 260170 280948 260176
rect 280804 253224 280856 253230
rect 280804 253166 280856 253172
rect 280896 209840 280948 209846
rect 280816 209788 280896 209794
rect 280816 209782 280948 209788
rect 280816 209778 280936 209782
rect 280804 209772 280936 209778
rect 280856 209766 280936 209772
rect 280804 209714 280856 209720
rect 280816 209683 280844 209714
rect 280988 200184 281040 200190
rect 280988 200126 281040 200132
rect 281000 200054 281028 200126
rect 280988 200048 281040 200054
rect 280988 199990 281040 199996
rect 280988 190868 281040 190874
rect 280988 190810 281040 190816
rect 281000 179382 281028 190810
rect 280988 179376 281040 179382
rect 280988 179318 281040 179324
rect 280986 172544 281042 172553
rect 280986 172479 281042 172488
rect 280804 171964 280856 171970
rect 280804 171906 280856 171912
rect 280816 162178 280844 171906
rect 280804 162172 280856 162178
rect 280804 162114 280856 162120
rect 281000 154601 281028 172479
rect 280986 154592 281042 154601
rect 280986 154527 281042 154536
rect 280804 152652 280856 152658
rect 280804 152594 280856 152600
rect 280816 152538 280844 152594
rect 62448 128336 62528 128364
rect 280724 152510 280844 152538
rect 62396 128318 62448 128324
rect 62394 128208 62450 128217
rect 62394 128143 62450 128152
rect 62408 116113 62436 128143
rect 280724 120136 280752 152510
rect 280804 152448 280856 152454
rect 280804 152390 280856 152396
rect 280816 125526 280844 152390
rect 280986 135280 281042 135289
rect 280986 135215 280988 135224
rect 281040 135215 281042 135224
rect 280988 135186 281040 135192
rect 280896 125724 280948 125730
rect 280896 125666 280948 125672
rect 280908 125594 280936 125666
rect 280896 125588 280948 125594
rect 280896 125530 280948 125536
rect 280804 125520 280856 125526
rect 280804 125462 280856 125468
rect 280804 120148 280856 120154
rect 280724 120108 280804 120136
rect 280804 120090 280856 120096
rect 280896 118652 280948 118658
rect 280896 118594 280948 118600
rect 62394 116104 62450 116113
rect 62394 116039 62450 116048
rect 280908 115954 280936 118594
rect 280908 115938 281028 115954
rect 280908 115932 281040 115938
rect 280908 115926 280988 115932
rect 280988 115874 281040 115880
rect 281000 115843 281028 115874
rect 280804 113960 280856 113966
rect 280724 113908 280804 113914
rect 280724 113902 280856 113908
rect 280724 113886 280844 113902
rect 62394 111480 62450 111489
rect 62394 111415 62450 111424
rect 62408 106321 62436 111415
rect 280724 106434 280752 113886
rect 280804 112396 280856 112402
rect 280804 112338 280856 112344
rect 280816 106554 280844 112338
rect 280804 106548 280856 106554
rect 280804 106490 280856 106496
rect 280724 106406 280844 106434
rect 62394 106312 62450 106321
rect 280816 106282 280844 106406
rect 280896 106344 280948 106350
rect 280896 106286 280948 106292
rect 62394 106247 62450 106256
rect 280804 106276 280856 106282
rect 280804 106218 280856 106224
rect 280908 106214 280936 106286
rect 280896 106208 280948 106214
rect 280896 106150 280948 106156
rect 62210 106040 62266 106049
rect 62210 105975 62266 105984
rect 62224 98297 62252 105975
rect 62316 98938 62528 98954
rect 62304 98932 62528 98938
rect 62356 98926 62528 98932
rect 62304 98874 62356 98880
rect 62210 98288 62266 98297
rect 62210 98223 62266 98232
rect 61382 98016 61438 98025
rect 61382 97951 61438 97960
rect 61396 97753 61424 97951
rect 61382 97744 61438 97753
rect 61382 97679 61438 97688
rect 62394 93800 62450 93809
rect 62394 93735 62450 93744
rect 62408 88641 62436 93735
rect 62394 88632 62450 88641
rect 62394 88567 62450 88576
rect 61382 86320 61438 86329
rect 61382 86255 61438 86264
rect 61292 43716 61344 43722
rect 61292 43658 61344 43664
rect 61396 38010 61424 86255
rect 62500 84946 62528 98926
rect 281092 96898 281120 262958
rect 281184 261594 281212 266970
rect 281262 266792 281318 266801
rect 281262 266727 281318 266736
rect 281172 261588 281224 261594
rect 281172 261530 281224 261536
rect 281276 260166 281304 266727
rect 281368 263566 281396 267242
rect 281356 263560 281408 263566
rect 281356 263502 281408 263508
rect 281264 260160 281316 260166
rect 281264 260102 281316 260108
rect 281170 219328 281226 219337
rect 281170 219263 281226 219272
rect 281184 209846 281212 219263
rect 281172 209840 281224 209846
rect 281172 209782 281224 209788
rect 281170 189680 281226 189689
rect 281170 189615 281226 189624
rect 281184 171970 281212 189615
rect 281448 179376 281500 179382
rect 281448 179318 281500 179324
rect 281172 171964 281224 171970
rect 281172 171906 281224 171912
rect 281460 166938 281488 179318
rect 281264 166932 281316 166938
rect 281264 166874 281316 166880
rect 281448 166932 281500 166938
rect 281448 166874 281500 166880
rect 281276 162330 281304 166874
rect 281184 162302 281304 162330
rect 281184 152658 281212 162302
rect 281264 162172 281316 162178
rect 281264 162114 281316 162120
rect 281172 152652 281224 152658
rect 281172 152594 281224 152600
rect 281276 152454 281304 162114
rect 281354 154592 281410 154601
rect 281354 154527 281410 154536
rect 281264 152448 281316 152454
rect 281264 152390 281316 152396
rect 281262 138544 281318 138553
rect 281262 138479 281318 138488
rect 281172 120148 281224 120154
rect 281172 120090 281224 120096
rect 281184 113966 281212 120090
rect 281172 113960 281224 113966
rect 281172 113902 281224 113908
rect 281172 106276 281224 106282
rect 281172 106218 281224 106224
rect 281080 96892 281132 96898
rect 281080 96834 281132 96840
rect 280988 96688 281040 96694
rect 280988 96630 281040 96636
rect 281080 96688 281132 96694
rect 281080 96630 281132 96636
rect 281000 96558 281028 96630
rect 280988 96552 281040 96558
rect 280988 96494 281040 96500
rect 280804 94648 280856 94654
rect 62224 84918 62528 84946
rect 280724 94596 280804 94602
rect 280724 94590 280856 94596
rect 280724 94574 280844 94590
rect 280724 84946 280752 94574
rect 280804 94512 280856 94518
rect 280804 94454 280856 94460
rect 280816 85066 280844 94454
rect 280988 89684 281040 89690
rect 280988 89626 281040 89632
rect 281000 86970 281028 89626
rect 280988 86964 281040 86970
rect 280988 86906 281040 86912
rect 280804 85060 280856 85066
rect 280804 85002 280856 85008
rect 280724 84930 280844 84946
rect 280724 84924 280856 84930
rect 280724 84918 280804 84924
rect 62224 77246 62252 84918
rect 280804 84866 280856 84872
rect 62394 81560 62450 81569
rect 62394 81495 62450 81504
rect 62302 79928 62358 79937
rect 62302 79863 62358 79872
rect 62212 77240 62264 77246
rect 62212 77182 62264 77188
rect 62210 70544 62266 70553
rect 62210 70479 62266 70488
rect 62224 60761 62252 70479
rect 62316 67833 62344 79863
rect 62302 67824 62358 67833
rect 62302 67759 62358 67768
rect 62304 67652 62356 67658
rect 62304 67594 62356 67600
rect 62210 60752 62266 60761
rect 62210 60687 62266 60696
rect 61474 58576 61530 58585
rect 61474 58511 61530 58520
rect 61488 43450 61516 58511
rect 62316 55842 62344 67594
rect 62132 55814 62344 55842
rect 62026 46336 62082 46345
rect 62026 46271 62082 46280
rect 62040 43654 62068 46271
rect 62028 43648 62080 43654
rect 62028 43590 62080 43596
rect 61476 43444 61528 43450
rect 61476 43386 61528 43392
rect 61384 38004 61436 38010
rect 61384 37946 61436 37952
rect 62132 35034 62160 55814
rect 62302 53952 62358 53961
rect 62302 53887 62358 53896
rect 62210 44976 62266 44985
rect 62210 44911 62266 44920
rect 62224 44334 62252 44911
rect 62212 44328 62264 44334
rect 62212 44270 62264 44276
rect 62316 35222 62344 53887
rect 62304 35216 62356 35222
rect 62304 35158 62356 35164
rect 62408 35154 62436 81495
rect 280908 77314 281028 77330
rect 280896 77308 281028 77314
rect 280948 77302 281028 77308
rect 280896 77250 280948 77256
rect 281000 77246 281028 77302
rect 280988 77240 281040 77246
rect 280988 77182 281040 77188
rect 280804 75336 280856 75342
rect 280724 75284 280804 75290
rect 280724 75278 280856 75284
rect 280724 75262 280844 75278
rect 280724 65498 280752 75262
rect 280804 75200 280856 75206
rect 280804 75142 280856 75148
rect 280816 67454 280844 75142
rect 280896 67720 280948 67726
rect 280896 67662 280948 67668
rect 280908 67590 280936 67662
rect 280896 67584 280948 67590
rect 280896 67526 280948 67532
rect 280804 67448 280856 67454
rect 280804 67390 280856 67396
rect 280724 65482 280844 65498
rect 280724 65476 280856 65482
rect 280724 65470 280804 65476
rect 280804 65418 280856 65424
rect 281092 60897 281120 96630
rect 281184 94654 281212 106218
rect 281172 94648 281224 94654
rect 281172 94590 281224 94596
rect 281170 84416 281226 84425
rect 281170 84351 281226 84360
rect 281078 60888 281134 60897
rect 281078 60823 281134 60832
rect 280988 60648 281040 60654
rect 280988 60590 281040 60596
rect 281000 51066 281028 60590
rect 281078 59664 281134 59673
rect 281078 59599 281134 59608
rect 280804 51060 280856 51066
rect 280804 51002 280856 51008
rect 280988 51060 281040 51066
rect 280988 51002 281040 51008
rect 280816 48278 280844 51002
rect 280896 48340 280948 48346
rect 280896 48282 280948 48288
rect 280804 48272 280856 48278
rect 280804 48214 280856 48220
rect 280908 44010 280936 48282
rect 280724 43982 280936 44010
rect 277032 43920 277084 43926
rect 277030 43888 277032 43897
rect 277084 43888 277086 43897
rect 144184 43852 144236 43858
rect 277030 43823 277086 43832
rect 144184 43794 144236 43800
rect 142066 43480 142122 43489
rect 142066 43415 142122 43424
rect 63512 40118 63540 43316
rect 64446 43302 64828 43330
rect 68494 43302 68968 43330
rect 64144 42968 64196 42974
rect 64144 42910 64196 42916
rect 63500 40112 63552 40118
rect 63500 40054 63552 40060
rect 62396 35148 62448 35154
rect 62396 35090 62448 35096
rect 62132 35006 62528 35034
rect 62396 34944 62448 34950
rect 62396 34886 62448 34892
rect 61200 25628 61252 25634
rect 61200 25570 61252 25576
rect 62408 19990 62436 34886
rect 62396 19984 62448 19990
rect 62396 19926 62448 19932
rect 61108 7812 61160 7818
rect 61108 7754 61160 7760
rect 57888 3936 57940 3942
rect 57888 3878 57940 3884
rect 57704 3664 57756 3670
rect 57704 3606 57756 3612
rect 62500 3398 62528 35006
rect 64156 3602 64184 42910
rect 64800 32502 64828 43302
rect 65524 40112 65576 40118
rect 65524 40054 65576 40060
rect 64788 32496 64840 32502
rect 64788 32438 64840 32444
rect 65536 7682 65564 40054
rect 68940 22982 68968 43302
rect 69400 40118 69428 43316
rect 70504 40118 70532 43316
rect 71438 43302 71636 43330
rect 69388 40112 69440 40118
rect 69388 40054 69440 40060
rect 70308 40112 70360 40118
rect 70308 40054 70360 40060
rect 70492 40112 70544 40118
rect 70492 40054 70544 40060
rect 70320 26926 70348 40054
rect 70308 26920 70360 26926
rect 70308 26862 70360 26868
rect 68928 22976 68980 22982
rect 68928 22918 68980 22924
rect 71608 14618 71636 43302
rect 71688 40112 71740 40118
rect 71688 40054 71740 40060
rect 71596 14612 71648 14618
rect 71596 14554 71648 14560
rect 65524 7676 65576 7682
rect 65524 7618 65576 7624
rect 71700 4826 71728 40054
rect 74368 39778 74396 43316
rect 79336 42809 79364 43316
rect 79322 42800 79378 42809
rect 79322 42735 79378 42744
rect 81360 39914 81388 43316
rect 81348 39908 81400 39914
rect 81348 39850 81400 39856
rect 82280 39846 82308 43316
rect 83200 40798 83228 43316
rect 83188 40792 83240 40798
rect 83188 40734 83240 40740
rect 84304 40118 84332 43316
rect 86328 42673 86356 43316
rect 86314 42664 86370 42673
rect 86314 42599 86370 42608
rect 87248 40866 87276 43316
rect 88168 41410 88196 43316
rect 88984 42084 89036 42090
rect 88984 42026 89036 42032
rect 88156 41404 88208 41410
rect 88156 41346 88208 41352
rect 88996 41274 89024 42026
rect 88984 41268 89036 41274
rect 88984 41210 89036 41216
rect 89272 41138 89300 43316
rect 89260 41132 89312 41138
rect 89260 41074 89312 41080
rect 87236 40860 87288 40866
rect 87236 40802 87288 40808
rect 91112 40118 91140 43316
rect 92230 43302 92428 43330
rect 84292 40112 84344 40118
rect 84292 40054 84344 40060
rect 85488 40112 85540 40118
rect 85488 40054 85540 40060
rect 91100 40112 91152 40118
rect 91100 40054 91152 40060
rect 92296 40112 92348 40118
rect 92296 40054 92348 40060
rect 82268 39840 82320 39846
rect 82268 39782 82320 39788
rect 74356 39772 74408 39778
rect 74356 39714 74408 39720
rect 85500 24410 85528 40054
rect 85488 24404 85540 24410
rect 85488 24346 85540 24352
rect 92308 10402 92336 40054
rect 92296 10396 92348 10402
rect 92296 10338 92348 10344
rect 92400 6322 92428 43302
rect 94240 42702 94268 43316
rect 94228 42696 94280 42702
rect 94228 42638 94280 42644
rect 95160 40050 95188 43316
rect 96080 40905 96108 43316
rect 96528 42288 96580 42294
rect 96528 42230 96580 42236
rect 96540 41410 96568 42230
rect 96528 41404 96580 41410
rect 96528 41346 96580 41352
rect 97184 41274 97212 43316
rect 97172 41268 97224 41274
rect 97172 41210 97224 41216
rect 96066 40896 96122 40905
rect 96066 40831 96122 40840
rect 95148 40044 95200 40050
rect 95148 39986 95200 39992
rect 99024 37330 99052 43316
rect 100128 41313 100156 43316
rect 100114 41304 100170 41313
rect 100114 41239 100170 41248
rect 101048 41177 101076 43316
rect 103086 43302 103468 43330
rect 101034 41168 101090 41177
rect 101034 41103 101090 41112
rect 99012 37324 99064 37330
rect 99012 37266 99064 37272
rect 99288 37324 99340 37330
rect 99288 37266 99340 37272
rect 99300 27606 99328 37266
rect 99288 27600 99340 27606
rect 99288 27542 99340 27548
rect 103440 17270 103468 43302
rect 103992 41138 104020 43316
rect 106016 41274 106044 43316
rect 106004 41268 106056 41274
rect 106004 41210 106056 41216
rect 103980 41132 104032 41138
rect 103980 41074 104032 41080
rect 106936 41070 106964 43316
rect 106924 41064 106976 41070
rect 106924 41006 106976 41012
rect 103428 17264 103480 17270
rect 103428 17206 103480 17212
rect 99196 9716 99248 9722
rect 99196 9658 99248 9664
rect 92388 6316 92440 6322
rect 92388 6258 92440 6264
rect 71688 4820 71740 4826
rect 71688 4762 71740 4768
rect 64144 3596 64196 3602
rect 64144 3538 64196 3544
rect 62488 3392 62540 3398
rect 57426 3360 57482 3369
rect 56508 3324 56560 3330
rect 62488 3334 62540 3340
rect 57426 3295 57482 3304
rect 56508 3266 56560 3272
rect 99208 3058 99236 9658
rect 108960 4894 108988 43316
rect 110984 40118 111012 43316
rect 111904 40730 111932 43316
rect 113022 43302 113128 43330
rect 111892 40724 111944 40730
rect 111892 40666 111944 40672
rect 110972 40112 111024 40118
rect 110972 40054 111024 40060
rect 111708 40112 111760 40118
rect 111708 40054 111760 40060
rect 111720 17338 111748 40054
rect 111708 17332 111760 17338
rect 111708 17274 111760 17280
rect 113100 9382 113128 43302
rect 114848 40118 114876 43316
rect 117990 43302 118648 43330
rect 115204 40792 115256 40798
rect 115204 40734 115256 40740
rect 114836 40112 114888 40118
rect 114836 40054 114888 40060
rect 113088 9376 113140 9382
rect 113088 9318 113140 9324
rect 108948 4888 109000 4894
rect 108948 4830 109000 4836
rect 115216 3534 115244 40734
rect 115848 40112 115900 40118
rect 115848 40054 115900 40060
rect 115860 15978 115888 40054
rect 118620 16114 118648 43302
rect 118896 40118 118924 43316
rect 119830 43302 120028 43330
rect 120934 43302 121408 43330
rect 118884 40112 118936 40118
rect 118884 40054 118936 40060
rect 119896 40112 119948 40118
rect 119896 40054 119948 40060
rect 119908 31278 119936 40054
rect 119896 31272 119948 31278
rect 119896 31214 119948 31220
rect 118608 16108 118660 16114
rect 118608 16050 118660 16056
rect 115848 15972 115900 15978
rect 115848 15914 115900 15920
rect 120000 6186 120028 43302
rect 121380 14482 121408 43302
rect 121458 42120 121514 42129
rect 121458 42055 121514 42064
rect 121472 41138 121500 42055
rect 121460 41132 121512 41138
rect 121460 41074 121512 41080
rect 121368 14476 121420 14482
rect 121368 14418 121420 14424
rect 122760 9450 122788 43316
rect 123878 43302 124168 43330
rect 124140 28558 124168 43302
rect 125888 40118 125916 43316
rect 126822 43302 126928 43330
rect 125876 40112 125928 40118
rect 125876 40054 125928 40060
rect 126796 40112 126848 40118
rect 126796 40054 126848 40060
rect 124128 28552 124180 28558
rect 124128 28494 124180 28500
rect 126808 25566 126836 40054
rect 126796 25560 126848 25566
rect 126796 25502 126848 25508
rect 122748 9444 122800 9450
rect 122748 9386 122800 9392
rect 126900 8974 126928 43302
rect 127728 41342 127756 43316
rect 128452 42152 128504 42158
rect 128452 42094 128504 42100
rect 128360 42084 128412 42090
rect 128360 42026 128412 42032
rect 127716 41336 127768 41342
rect 127716 41278 127768 41284
rect 128372 41274 128400 42026
rect 128360 41268 128412 41274
rect 128360 41210 128412 41216
rect 128268 29708 128320 29714
rect 128268 29650 128320 29656
rect 126888 8968 126940 8974
rect 126888 8910 126940 8916
rect 119988 6180 120040 6186
rect 119988 6122 120040 6128
rect 126610 3904 126666 3913
rect 126610 3839 126666 3848
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 122748 3392 122800 3398
rect 122748 3334 122800 3340
rect 122760 3058 122788 3334
rect 99196 3052 99248 3058
rect 99196 2994 99248 3000
rect 122748 3052 122800 3058
rect 122748 2994 122800 3000
rect 126624 480 126652 3839
rect 128280 3330 128308 29650
rect 128464 3466 128492 42094
rect 128832 41002 128860 43316
rect 128820 40996 128872 41002
rect 128820 40938 128872 40944
rect 129648 40996 129700 41002
rect 129648 40938 129700 40944
rect 129660 18902 129688 40938
rect 129752 40118 129780 43316
rect 130686 43302 130976 43330
rect 131790 43302 132448 43330
rect 129740 40112 129792 40118
rect 129740 40054 129792 40060
rect 130948 22914 130976 43302
rect 131028 40112 131080 40118
rect 131028 40054 131080 40060
rect 130936 22908 130988 22914
rect 130936 22850 130988 22856
rect 131040 21418 131068 40054
rect 131028 21412 131080 21418
rect 131028 21354 131080 21360
rect 129648 18896 129700 18902
rect 129648 18838 129700 18844
rect 131396 11960 131448 11966
rect 131396 11902 131448 11908
rect 128452 3460 128504 3466
rect 128452 3402 128504 3408
rect 129004 3460 129056 3466
rect 129004 3402 129056 3408
rect 127808 3324 127860 3330
rect 127808 3266 127860 3272
rect 128268 3324 128320 3330
rect 128268 3266 128320 3272
rect 127820 480 127848 3266
rect 129016 480 129044 3402
rect 130200 3188 130252 3194
rect 130200 3130 130252 3136
rect 130212 480 130240 3130
rect 131408 480 131436 11902
rect 132420 5098 132448 43302
rect 132696 40118 132724 43316
rect 134734 43302 135116 43330
rect 132684 40112 132736 40118
rect 132684 40054 132736 40060
rect 133788 40112 133840 40118
rect 133788 40054 133840 40060
rect 133604 11892 133656 11898
rect 133604 11834 133656 11840
rect 132408 5092 132460 5098
rect 132408 5034 132460 5040
rect 132592 3052 132644 3058
rect 132592 2994 132644 3000
rect 132604 480 132632 2994
rect 133616 2802 133644 11834
rect 133800 6390 133828 40054
rect 135088 24138 135116 43302
rect 135640 40118 135668 43316
rect 136744 40118 136772 43316
rect 138598 43302 139256 43330
rect 137008 41336 137060 41342
rect 137008 41278 137060 41284
rect 135628 40112 135680 40118
rect 135628 40054 135680 40060
rect 136456 40112 136508 40118
rect 136456 40054 136508 40060
rect 136732 40112 136784 40118
rect 136732 40054 136784 40060
rect 135168 38684 135220 38690
rect 135168 38626 135220 38632
rect 135180 38554 135208 38626
rect 135168 38548 135220 38554
rect 135168 38490 135220 38496
rect 135168 29028 135220 29034
rect 135168 28970 135220 28976
rect 135076 24132 135128 24138
rect 135076 24074 135128 24080
rect 135180 19650 135208 28970
rect 135168 19644 135220 19650
rect 135168 19586 135220 19592
rect 135168 19372 135220 19378
rect 135168 19314 135220 19320
rect 135180 19242 135208 19314
rect 135168 19236 135220 19242
rect 135168 19178 135220 19184
rect 136468 12034 136496 40054
rect 136546 39264 136602 39273
rect 136546 39199 136602 39208
rect 136456 12028 136508 12034
rect 136456 11970 136508 11976
rect 134892 9716 134944 9722
rect 134892 9658 134944 9664
rect 133788 6384 133840 6390
rect 133788 6326 133840 6332
rect 133616 2774 133828 2802
rect 133800 480 133828 2774
rect 134904 480 134932 9658
rect 136560 3466 136588 39199
rect 137020 38622 137048 41278
rect 137928 40112 137980 40118
rect 137928 40054 137980 40060
rect 137008 38616 137060 38622
rect 137008 38558 137060 38564
rect 137100 29028 137152 29034
rect 137100 28970 137152 28976
rect 137112 22114 137140 28970
rect 136928 22086 137140 22114
rect 136928 12458 136956 22086
rect 137940 13122 137968 40054
rect 139228 21554 139256 43302
rect 139688 41070 139716 43316
rect 140622 43302 140728 43330
rect 141726 43302 142016 43330
rect 139676 41064 139728 41070
rect 139676 41006 139728 41012
rect 139306 29880 139362 29889
rect 139306 29815 139362 29824
rect 139216 21548 139268 21554
rect 139216 21490 139268 21496
rect 137928 13116 137980 13122
rect 137928 13058 137980 13064
rect 136744 12430 136956 12458
rect 136744 3466 136772 12430
rect 139320 3466 139348 29815
rect 140700 14550 140728 43302
rect 141988 28354 142016 43302
rect 141976 28348 142028 28354
rect 141976 28290 142028 28296
rect 140688 14544 140740 14550
rect 140688 14486 140740 14492
rect 142080 3466 142108 43415
rect 142632 40118 142660 43316
rect 143552 41206 143580 43316
rect 143540 41200 143592 41206
rect 143540 41142 143592 41148
rect 142620 40112 142672 40118
rect 142620 40054 142672 40060
rect 143448 40112 143500 40118
rect 143448 40054 143500 40060
rect 143356 18828 143408 18834
rect 143356 18770 143408 18776
rect 143368 3482 143396 18770
rect 143460 5030 143488 40054
rect 143448 5024 143500 5030
rect 143448 4966 143500 4972
rect 136088 3460 136140 3466
rect 136088 3402 136140 3408
rect 136548 3460 136600 3466
rect 136548 3402 136600 3408
rect 136732 3460 136784 3466
rect 136732 3402 136784 3408
rect 137284 3460 137336 3466
rect 137284 3402 137336 3408
rect 138480 3460 138532 3466
rect 138480 3402 138532 3408
rect 139308 3460 139360 3466
rect 139308 3402 139360 3408
rect 140872 3460 140924 3466
rect 140872 3402 140924 3408
rect 142068 3460 142120 3466
rect 142068 3402 142120 3408
rect 143276 3454 143396 3482
rect 144196 3466 144224 43794
rect 187700 43716 187752 43722
rect 187700 43658 187752 43664
rect 211068 43716 211120 43722
rect 211068 43658 211120 43664
rect 151004 43438 151478 43466
rect 144670 43302 144868 43330
rect 145590 43302 146248 43330
rect 144840 22778 144868 43302
rect 146220 31142 146248 43302
rect 146496 42566 146524 43316
rect 146588 43302 147614 43330
rect 148534 43302 148916 43330
rect 146484 42560 146536 42566
rect 146484 42502 146536 42508
rect 146588 33794 146616 43302
rect 146576 33788 146628 33794
rect 146576 33730 146628 33736
rect 146208 31136 146260 31142
rect 146208 31078 146260 31084
rect 146668 29028 146720 29034
rect 146668 28970 146720 28976
rect 146298 28248 146354 28257
rect 146298 28183 146354 28192
rect 144828 22772 144880 22778
rect 144828 22714 144880 22720
rect 144460 6724 144512 6730
rect 144460 6666 144512 6672
rect 144184 3460 144236 3466
rect 136100 480 136128 3402
rect 137296 480 137324 3402
rect 138492 480 138520 3402
rect 139674 3224 139730 3233
rect 139674 3159 139730 3168
rect 139688 480 139716 3159
rect 140884 480 140912 3402
rect 142068 3256 142120 3262
rect 142068 3198 142120 3204
rect 142080 480 142108 3198
rect 143276 480 143304 3454
rect 144184 3402 144236 3408
rect 144472 480 144500 6666
rect 145656 3460 145708 3466
rect 145656 3402 145708 3408
rect 145668 480 145696 3402
rect 146312 3346 146340 28183
rect 146680 22098 146708 28970
rect 148888 24342 148916 43302
rect 149624 40118 149652 43316
rect 151004 40338 151032 43438
rect 152582 43302 153056 43330
rect 150820 40310 151032 40338
rect 149612 40112 149664 40118
rect 149612 40054 149664 40060
rect 150348 40112 150400 40118
rect 150348 40054 150400 40060
rect 149060 37324 149112 37330
rect 149060 37266 149112 37272
rect 149072 27606 149100 37266
rect 149060 27600 149112 27606
rect 149060 27542 149112 27548
rect 148968 25696 149020 25702
rect 148968 25638 149020 25644
rect 148876 24336 148928 24342
rect 148876 24278 148928 24284
rect 146668 22092 146720 22098
rect 146668 22034 146720 22040
rect 148980 3466 149008 25638
rect 149060 18012 149112 18018
rect 149060 17954 149112 17960
rect 149072 12510 149100 17954
rect 149060 12504 149112 12510
rect 149060 12446 149112 12452
rect 149244 12300 149296 12306
rect 149244 12242 149296 12248
rect 148048 3460 148100 3466
rect 148048 3402 148100 3408
rect 148968 3460 149020 3466
rect 148968 3402 149020 3408
rect 146312 3318 146892 3346
rect 146864 480 146892 3318
rect 148060 480 148088 3402
rect 149256 480 149284 12242
rect 150360 3398 150388 40054
rect 150820 29073 150848 40310
rect 150622 29064 150678 29073
rect 150622 28999 150678 29008
rect 150806 29064 150862 29073
rect 150806 28999 150862 29008
rect 150636 27606 150664 28999
rect 153028 28490 153056 43302
rect 153106 42256 153162 42265
rect 153106 42191 153162 42200
rect 153016 28484 153068 28490
rect 153016 28426 153068 28432
rect 150624 27600 150676 27606
rect 150624 27542 150676 27548
rect 150716 11688 150768 11694
rect 150716 11630 150768 11636
rect 150728 3466 150756 11630
rect 150716 3460 150768 3466
rect 150716 3402 150768 3408
rect 151544 3460 151596 3466
rect 151544 3402 151596 3408
rect 150348 3392 150400 3398
rect 150348 3334 150400 3340
rect 150440 3324 150492 3330
rect 150440 3266 150492 3272
rect 150452 480 150480 3266
rect 151556 480 151584 3402
rect 153120 2854 153148 42191
rect 153488 41002 153516 43316
rect 155526 43302 155816 43330
rect 154488 42220 154540 42226
rect 154488 42162 154540 42168
rect 153476 40996 153528 41002
rect 153476 40938 153528 40944
rect 154500 3466 154528 42162
rect 155788 10470 155816 43302
rect 157248 42356 157300 42362
rect 157248 42298 157300 42304
rect 155868 42288 155920 42294
rect 155868 42230 155920 42236
rect 155776 10464 155828 10470
rect 155776 10406 155828 10412
rect 155880 3466 155908 42230
rect 153936 3460 153988 3466
rect 153936 3402 153988 3408
rect 154488 3460 154540 3466
rect 154488 3402 154540 3408
rect 155132 3460 155184 3466
rect 155132 3402 155184 3408
rect 155868 3460 155920 3466
rect 155868 3402 155920 3408
rect 153108 2848 153160 2854
rect 153108 2790 153160 2796
rect 152740 604 152792 610
rect 152740 546 152792 552
rect 152752 480 152780 546
rect 153948 480 153976 3402
rect 155144 480 155172 3402
rect 157260 3398 157288 42298
rect 157536 40118 157564 43316
rect 158456 42537 158484 43316
rect 160480 42634 160508 43316
rect 160468 42628 160520 42634
rect 160468 42570 160520 42576
rect 158442 42528 158498 42537
rect 158442 42463 158498 42472
rect 161400 42401 161428 43316
rect 162334 43302 162808 43330
rect 161386 42392 161442 42401
rect 161386 42327 161442 42336
rect 158628 41132 158680 41138
rect 158628 41074 158680 41080
rect 157524 40112 157576 40118
rect 157524 40054 157576 40060
rect 158536 40112 158588 40118
rect 158536 40054 158588 40060
rect 158548 28286 158576 40054
rect 158536 28280 158588 28286
rect 158536 28222 158588 28228
rect 158640 3398 158668 41074
rect 162676 21480 162728 21486
rect 162676 21422 162728 21428
rect 160006 16008 160062 16017
rect 160006 15943 160062 15952
rect 159916 7948 159968 7954
rect 159916 7890 159968 7896
rect 156328 3392 156380 3398
rect 156328 3334 156380 3340
rect 157248 3392 157300 3398
rect 157248 3334 157300 3340
rect 157524 3392 157576 3398
rect 157524 3334 157576 3340
rect 158628 3392 158680 3398
rect 158628 3334 158680 3340
rect 158720 3392 158772 3398
rect 158720 3334 158772 3340
rect 156340 480 156368 3334
rect 157536 480 157564 3334
rect 158732 480 158760 3334
rect 159928 480 159956 7890
rect 160020 3398 160048 15943
rect 161112 4140 161164 4146
rect 161112 4082 161164 4088
rect 160008 3392 160060 3398
rect 160008 3334 160060 3340
rect 161124 480 161152 4082
rect 162688 3482 162716 21422
rect 162780 9586 162808 43302
rect 163424 40118 163452 43316
rect 164344 40798 164372 43316
rect 164332 40792 164384 40798
rect 164332 40734 164384 40740
rect 167288 40118 167316 43316
rect 168288 42424 168340 42430
rect 168288 42366 168340 42372
rect 163412 40112 163464 40118
rect 163412 40054 163464 40060
rect 164148 40112 164200 40118
rect 164148 40054 164200 40060
rect 167276 40112 167328 40118
rect 167276 40054 167328 40060
rect 168196 40112 168248 40118
rect 168196 40054 168248 40060
rect 164160 33182 164188 40054
rect 164148 33176 164200 33182
rect 164148 33118 164200 33124
rect 162860 19984 162912 19990
rect 162860 19926 162912 19932
rect 162768 9580 162820 9586
rect 162768 9522 162820 9528
rect 162320 3454 162716 3482
rect 162872 3482 162900 19926
rect 168208 17542 168236 40054
rect 168196 17536 168248 17542
rect 168196 17478 168248 17484
rect 166908 12096 166960 12102
rect 166908 12038 166960 12044
rect 164700 4072 164752 4078
rect 164700 4014 164752 4020
rect 162872 3454 163544 3482
rect 162320 480 162348 3454
rect 163516 480 163544 3454
rect 164712 480 164740 4014
rect 166920 2990 166948 12038
rect 167000 12028 167052 12034
rect 167000 11970 167052 11976
rect 167012 3482 167040 11970
rect 168300 3482 168328 42366
rect 168392 41177 168420 43316
rect 169326 43302 169708 43330
rect 168378 41168 168434 41177
rect 168378 41103 168434 41112
rect 168380 33176 168432 33182
rect 168380 33118 168432 33124
rect 167012 3454 167132 3482
rect 165896 2984 165948 2990
rect 165896 2926 165948 2932
rect 166908 2984 166960 2990
rect 166908 2926 166960 2932
rect 165908 480 165936 2926
rect 167104 480 167132 3454
rect 168208 3454 168328 3482
rect 168392 3482 168420 33118
rect 169680 9654 169708 43302
rect 170232 40118 170260 43316
rect 171336 40118 171364 43316
rect 172270 43302 172468 43330
rect 173374 43302 173848 43330
rect 170220 40112 170272 40118
rect 170220 40054 170272 40060
rect 171048 40112 171100 40118
rect 171048 40054 171100 40060
rect 171324 40112 171376 40118
rect 171324 40054 171376 40060
rect 172336 40112 172388 40118
rect 172336 40054 172388 40060
rect 170956 25764 171008 25770
rect 170956 25706 171008 25712
rect 169668 9648 169720 9654
rect 169668 9590 169720 9596
rect 170968 3482 170996 25706
rect 171060 10538 171088 40054
rect 172348 33794 172376 40054
rect 172336 33788 172388 33794
rect 172336 33730 172388 33736
rect 172440 10674 172468 43302
rect 173820 20618 173848 43302
rect 174280 40118 174308 43316
rect 178144 40118 178172 43316
rect 179156 43302 179262 43330
rect 180182 43302 180748 43330
rect 174268 40112 174320 40118
rect 174268 40054 174320 40060
rect 175188 40112 175240 40118
rect 175188 40054 175240 40060
rect 178132 40112 178184 40118
rect 178132 40054 178184 40060
rect 173820 20590 173940 20618
rect 172428 10668 172480 10674
rect 172428 10610 172480 10616
rect 171048 10532 171100 10538
rect 171048 10474 171100 10480
rect 172978 6896 173034 6905
rect 172978 6831 173034 6840
rect 171782 3768 171838 3777
rect 171782 3703 171838 3712
rect 168392 3454 169432 3482
rect 168208 480 168236 3454
rect 169404 480 169432 3454
rect 170600 3454 170996 3482
rect 170600 480 170628 3454
rect 171796 480 171824 3703
rect 172992 480 173020 6831
rect 173912 3482 173940 20590
rect 175200 18698 175228 40054
rect 179156 32570 179184 43302
rect 179236 40112 179288 40118
rect 179236 40054 179288 40060
rect 179144 32564 179196 32570
rect 179144 32506 179196 32512
rect 176568 23044 176620 23050
rect 176568 22986 176620 22992
rect 175188 18692 175240 18698
rect 175188 18634 175240 18640
rect 176476 4004 176528 4010
rect 176476 3946 176528 3952
rect 173912 3454 174216 3482
rect 174188 480 174216 3454
rect 175372 3392 175424 3398
rect 175372 3334 175424 3340
rect 175384 480 175412 3334
rect 176488 3210 176516 3946
rect 176580 3398 176608 22986
rect 179248 19990 179276 40054
rect 179328 36712 179380 36718
rect 179328 36654 179380 36660
rect 179236 19984 179288 19990
rect 179236 19926 179288 19932
rect 177764 6656 177816 6662
rect 177764 6598 177816 6604
rect 176568 3392 176620 3398
rect 176568 3334 176620 3340
rect 176488 3182 176608 3210
rect 176580 480 176608 3182
rect 177776 480 177804 6598
rect 179340 3482 179368 36654
rect 180720 9246 180748 43302
rect 181272 41274 181300 43316
rect 181260 41268 181312 41274
rect 181260 41210 181312 41216
rect 182088 41268 182140 41274
rect 182088 41210 182140 41216
rect 182100 18766 182128 41210
rect 182192 40118 182220 43316
rect 183126 43302 183508 43330
rect 184230 43302 184888 43330
rect 182180 40112 182232 40118
rect 182180 40054 182232 40060
rect 183376 40112 183428 40118
rect 183376 40054 183428 40060
rect 182088 18760 182140 18766
rect 182088 18702 182140 18708
rect 182088 13796 182140 13802
rect 182088 13738 182140 13744
rect 180708 9240 180760 9246
rect 180708 9182 180760 9188
rect 180156 5228 180208 5234
rect 180156 5170 180208 5176
rect 178972 3454 179368 3482
rect 178972 480 179000 3454
rect 180168 480 180196 5170
rect 182100 3398 182128 13738
rect 183388 12034 183416 40054
rect 183376 12028 183428 12034
rect 183376 11970 183428 11976
rect 182548 6656 182600 6662
rect 182548 6598 182600 6604
rect 181352 3392 181404 3398
rect 181352 3334 181404 3340
rect 182088 3392 182140 3398
rect 182088 3334 182140 3340
rect 181364 480 181392 3334
rect 182560 480 182588 6598
rect 183480 5166 183508 43302
rect 183558 30968 183614 30977
rect 183558 30903 183614 30912
rect 183468 5160 183520 5166
rect 183468 5102 183520 5108
rect 183572 3398 183600 30903
rect 184860 7886 184888 43302
rect 185136 42634 185164 43316
rect 185596 43302 186070 43330
rect 187174 43302 187648 43330
rect 185124 42628 185176 42634
rect 185124 42570 185176 42576
rect 185596 31906 185624 43302
rect 186320 39432 186372 39438
rect 186320 39374 186372 39380
rect 185320 31878 185624 31906
rect 185320 31770 185348 31878
rect 185136 31742 185348 31770
rect 185136 13802 185164 31742
rect 185124 13796 185176 13802
rect 185124 13738 185176 13744
rect 184848 7880 184900 7886
rect 184848 7822 184900 7828
rect 183744 4004 183796 4010
rect 183744 3946 183796 3952
rect 183560 3392 183612 3398
rect 183560 3334 183612 3340
rect 183756 480 183784 3946
rect 186044 3936 186096 3942
rect 186044 3878 186096 3884
rect 184848 3392 184900 3398
rect 184848 3334 184900 3340
rect 184860 480 184888 3334
rect 186056 480 186084 3878
rect 186332 610 186360 39374
rect 187620 9518 187648 43302
rect 187608 9512 187660 9518
rect 187608 9454 187660 9460
rect 187712 610 187740 43658
rect 189184 40118 189212 43316
rect 190104 41993 190132 43316
rect 191024 42566 191052 43316
rect 193062 43302 193168 43330
rect 191012 42560 191064 42566
rect 191012 42502 191064 42508
rect 190090 41984 190146 41993
rect 190090 41919 190146 41928
rect 189172 40112 189224 40118
rect 189172 40054 189224 40060
rect 190368 40112 190420 40118
rect 190368 40054 190420 40060
rect 190380 13190 190408 40054
rect 190368 13184 190420 13190
rect 190368 13126 190420 13132
rect 193140 10606 193168 43302
rect 195072 42498 195100 43316
rect 195060 42492 195112 42498
rect 195060 42434 195112 42440
rect 195992 40118 196020 43316
rect 197110 43302 197308 43330
rect 195980 40112 196032 40118
rect 195980 40054 196032 40060
rect 197176 40112 197228 40118
rect 197176 40054 197228 40060
rect 194506 39400 194562 39409
rect 194506 39335 194562 39344
rect 193220 38004 193272 38010
rect 193220 37946 193272 37952
rect 193128 10600 193180 10606
rect 193128 10542 193180 10548
rect 189632 8832 189684 8838
rect 189632 8774 189684 8780
rect 186320 604 186372 610
rect 186320 546 186372 552
rect 187240 604 187292 610
rect 187240 546 187292 552
rect 187700 604 187752 610
rect 187700 546 187752 552
rect 188436 604 188488 610
rect 188436 546 188488 552
rect 187252 480 187280 546
rect 188448 480 188476 546
rect 189644 480 189672 8774
rect 192024 6792 192076 6798
rect 192024 6734 192076 6740
rect 190828 3868 190880 3874
rect 190828 3810 190880 3816
rect 190840 480 190868 3810
rect 192036 480 192064 6734
rect 193232 2922 193260 37946
rect 193220 2916 193272 2922
rect 193220 2858 193272 2864
rect 194416 2916 194468 2922
rect 194416 2858 194468 2864
rect 193220 2780 193272 2786
rect 193220 2722 193272 2728
rect 193232 480 193260 2722
rect 194428 480 194456 2858
rect 194520 2854 194548 39335
rect 197188 15910 197216 40054
rect 197176 15904 197228 15910
rect 197176 15846 197228 15852
rect 196808 8900 196860 8906
rect 196808 8842 196860 8848
rect 195612 6452 195664 6458
rect 195612 6394 195664 6400
rect 194508 2848 194560 2854
rect 194508 2790 194560 2796
rect 195624 480 195652 6394
rect 196820 480 196848 8842
rect 197280 4962 197308 43302
rect 198016 41206 198044 43316
rect 198752 43302 198950 43330
rect 198004 41200 198056 41206
rect 198004 41142 198056 41148
rect 198752 5234 198780 43302
rect 200040 42906 200068 43316
rect 200028 42900 200080 42906
rect 200028 42842 200080 42848
rect 202984 40118 203012 43316
rect 203918 43302 204208 43330
rect 205022 43302 205588 43330
rect 202972 40112 203024 40118
rect 202972 40054 203024 40060
rect 204076 40112 204128 40118
rect 204076 40054 204128 40060
rect 202788 38004 202840 38010
rect 202788 37946 202840 37952
rect 198740 5228 198792 5234
rect 198740 5170 198792 5176
rect 201500 5092 201552 5098
rect 201500 5034 201552 5040
rect 197268 4956 197320 4962
rect 197268 4898 197320 4904
rect 199200 3936 199252 3942
rect 199200 3878 199252 3884
rect 198004 3664 198056 3670
rect 198004 3606 198056 3612
rect 198016 480 198044 3606
rect 199212 480 199240 3878
rect 200394 3632 200450 3641
rect 200394 3567 200450 3576
rect 200408 480 200436 3567
rect 201512 480 201540 5034
rect 202800 3482 202828 37946
rect 203984 20052 204036 20058
rect 203984 19994 204036 20000
rect 203996 3482 204024 19994
rect 204088 17474 204116 40054
rect 204076 17468 204128 17474
rect 204076 17410 204128 17416
rect 204180 7614 204208 43302
rect 204904 41200 204956 41206
rect 204904 41142 204956 41148
rect 204168 7608 204220 7614
rect 204168 7550 204220 7556
rect 204916 3670 204944 41142
rect 205560 10742 205588 43302
rect 205928 42537 205956 43316
rect 207966 43302 208256 43330
rect 205914 42528 205970 42537
rect 205914 42463 205970 42472
rect 205548 10736 205600 10742
rect 205548 10678 205600 10684
rect 208228 8022 208256 43302
rect 208308 41200 208360 41206
rect 208308 41142 208360 41148
rect 208216 8016 208268 8022
rect 208216 7958 208268 7964
rect 205088 4072 205140 4078
rect 205088 4014 205140 4020
rect 204904 3664 204956 3670
rect 204904 3606 204956 3612
rect 202708 3454 202828 3482
rect 203904 3454 204024 3482
rect 202708 480 202736 3454
rect 203904 480 203932 3454
rect 205100 480 205128 4014
rect 206284 3596 206336 3602
rect 206284 3538 206336 3544
rect 206296 480 206324 3538
rect 208320 3058 208348 41142
rect 209792 40118 209820 43316
rect 210896 41274 210924 43316
rect 210884 41268 210936 41274
rect 210884 41210 210936 41216
rect 209780 40112 209832 40118
rect 209780 40054 209832 40060
rect 210976 40112 211028 40118
rect 210976 40054 211028 40060
rect 210988 14686 211016 40054
rect 210976 14680 211028 14686
rect 210976 14622 211028 14628
rect 209870 6080 209926 6089
rect 209870 6015 209926 6024
rect 208676 5092 208728 5098
rect 208676 5034 208728 5040
rect 207480 3052 207532 3058
rect 207480 2994 207532 3000
rect 208308 3052 208360 3058
rect 208308 2994 208360 3000
rect 207492 480 207520 2994
rect 208688 480 208716 5034
rect 209884 480 209912 6015
rect 211080 480 211108 43658
rect 223856 43648 223908 43654
rect 223856 43590 223908 43596
rect 211816 41206 211844 43316
rect 211804 41200 211856 41206
rect 211804 41142 211856 41148
rect 212920 40118 212948 43316
rect 212908 40112 212960 40118
rect 212908 40054 212960 40060
rect 213736 40112 213788 40118
rect 213736 40054 213788 40060
rect 213748 32434 213776 40054
rect 213736 32428 213788 32434
rect 213736 32370 213788 32376
rect 213840 7750 213868 43316
rect 214774 43302 215248 43330
rect 215220 24274 215248 43302
rect 215864 40118 215892 43316
rect 216784 41410 216812 43316
rect 216772 41404 216824 41410
rect 216772 41346 216824 41352
rect 215852 40112 215904 40118
rect 215852 40054 215904 40060
rect 216588 40112 216640 40118
rect 216588 40054 216640 40060
rect 215208 24268 215260 24274
rect 215208 24210 215260 24216
rect 214656 8016 214708 8022
rect 214656 7958 214708 7964
rect 213828 7744 213880 7750
rect 213828 7686 213880 7692
rect 212264 6860 212316 6866
rect 212264 6802 212316 6808
rect 212276 480 212304 6802
rect 213460 6248 213512 6254
rect 213460 6190 213512 6196
rect 213472 480 213500 6190
rect 214668 480 214696 7958
rect 215852 5160 215904 5166
rect 215852 5102 215904 5108
rect 215864 480 215892 5102
rect 216600 3602 216628 40054
rect 219728 39710 219756 43316
rect 220832 40118 220860 43316
rect 221752 41041 221780 43316
rect 223684 43302 223790 43330
rect 221738 41032 221794 41041
rect 221738 40967 221794 40976
rect 220820 40112 220872 40118
rect 220820 40054 220872 40060
rect 222108 40112 222160 40118
rect 222108 40054 222160 40060
rect 219716 39704 219768 39710
rect 219716 39646 219768 39652
rect 219348 33924 219400 33930
rect 219348 33866 219400 33872
rect 218152 8764 218204 8770
rect 218152 8706 218204 8712
rect 217048 3868 217100 3874
rect 217048 3810 217100 3816
rect 216588 3596 216640 3602
rect 216588 3538 216640 3544
rect 217060 480 217088 3810
rect 218164 480 218192 8706
rect 219360 480 219388 33866
rect 220728 24472 220780 24478
rect 220728 24414 220780 24420
rect 220740 3482 220768 24414
rect 221740 7812 221792 7818
rect 221740 7754 221792 7760
rect 220556 3454 220768 3482
rect 220556 480 220584 3454
rect 221752 480 221780 7754
rect 222120 5166 222148 40054
rect 223212 32496 223264 32502
rect 223212 32438 223264 32444
rect 223224 30326 223252 32438
rect 223212 30320 223264 30326
rect 223212 30262 223264 30268
rect 223684 6730 223712 43302
rect 223672 6724 223724 6730
rect 223672 6666 223724 6672
rect 222108 5160 222160 5166
rect 222108 5102 222160 5108
rect 222936 3800 222988 3806
rect 222936 3742 222988 3748
rect 222948 480 222976 3742
rect 223868 3482 223896 43590
rect 227720 43580 227772 43586
rect 227720 43522 227772 43528
rect 224710 43302 224908 43330
rect 225630 43302 226288 43330
rect 224880 7818 224908 43302
rect 225328 9240 225380 9246
rect 225328 9182 225380 9188
rect 224868 7812 224920 7818
rect 224868 7754 224920 7760
rect 223868 3454 224172 3482
rect 224144 480 224172 3454
rect 225340 480 225368 9182
rect 226260 6458 226288 43302
rect 226340 31136 226392 31142
rect 226340 31078 226392 31084
rect 226248 6452 226300 6458
rect 226248 6394 226300 6400
rect 226352 3482 226380 31078
rect 226352 3454 226564 3482
rect 226536 480 226564 3454
rect 227732 480 227760 43522
rect 280724 43466 280752 43982
rect 237668 43438 238510 43466
rect 280632 43438 280752 43466
rect 229664 41274 229692 43316
rect 229652 41268 229704 41274
rect 229652 41210 229704 41216
rect 230584 40118 230612 43316
rect 233528 42838 233556 43316
rect 233516 42832 233568 42838
rect 233516 42774 233568 42780
rect 234632 41138 234660 43316
rect 234620 41132 234672 41138
rect 234620 41074 234672 41080
rect 235552 40934 235580 43316
rect 237392 43302 237590 43330
rect 235540 40928 235592 40934
rect 235540 40870 235592 40876
rect 230572 40112 230624 40118
rect 230572 40054 230624 40060
rect 231768 40112 231820 40118
rect 231768 40054 231820 40060
rect 231780 28626 231808 40054
rect 231768 28620 231820 28626
rect 231768 28562 231820 28568
rect 234620 28552 234672 28558
rect 234620 28494 234672 28500
rect 233240 24404 233292 24410
rect 233240 24346 233292 24352
rect 231768 16176 231820 16182
rect 231768 16118 231820 16124
rect 228916 8968 228968 8974
rect 228916 8910 228968 8916
rect 228928 480 228956 8910
rect 230112 5160 230164 5166
rect 230112 5102 230164 5108
rect 230124 480 230152 5102
rect 231780 3398 231808 16118
rect 232502 3632 232558 3641
rect 232502 3567 232558 3576
rect 231308 3392 231360 3398
rect 231308 3334 231360 3340
rect 231768 3392 231820 3398
rect 231768 3334 231820 3340
rect 231320 480 231348 3334
rect 232516 480 232544 3567
rect 233252 3482 233280 24346
rect 234632 14498 234660 28494
rect 236000 25628 236052 25634
rect 236000 25570 236052 25576
rect 234540 14470 234660 14498
rect 234540 9722 234568 14470
rect 234528 9716 234580 9722
rect 234528 9658 234580 9664
rect 234804 9716 234856 9722
rect 234804 9658 234856 9664
rect 233252 3454 233740 3482
rect 233712 480 233740 3454
rect 234816 480 234844 9658
rect 236012 480 236040 25570
rect 236092 14612 236144 14618
rect 236092 14554 236144 14560
rect 236104 610 236132 14554
rect 237392 8770 237420 43302
rect 237668 31890 237696 43438
rect 239404 41268 239456 41274
rect 239404 41210 239456 41216
rect 237656 31884 237708 31890
rect 237656 31826 237708 31832
rect 237656 31748 237708 31754
rect 237656 31690 237708 31696
rect 237668 22114 237696 31690
rect 237668 22086 237788 22114
rect 237564 18896 237616 18902
rect 237564 18838 237616 18844
rect 237472 12504 237524 12510
rect 237472 12446 237524 12452
rect 237484 11898 237512 12446
rect 237472 11892 237524 11898
rect 237472 11834 237524 11840
rect 237380 8764 237432 8770
rect 237380 8706 237432 8712
rect 237576 610 237604 18838
rect 237760 12510 237788 22086
rect 237748 12504 237800 12510
rect 237748 12446 237800 12452
rect 239416 9246 239444 41210
rect 239600 41206 239628 43316
rect 239588 41200 239640 41206
rect 239588 41142 239640 41148
rect 240520 40254 240548 43316
rect 241348 43302 241454 43330
rect 241532 43302 242558 43330
rect 240508 40248 240560 40254
rect 240508 40190 240560 40196
rect 241244 40248 241296 40254
rect 241244 40190 241296 40196
rect 241256 25634 241284 40190
rect 241244 25628 241296 25634
rect 241244 25570 241296 25576
rect 240048 14612 240100 14618
rect 240048 14554 240100 14560
rect 239404 9240 239456 9246
rect 239404 9182 239456 9188
rect 240060 4146 240088 14554
rect 241348 6254 241376 43302
rect 241428 38072 241480 38078
rect 241428 38014 241480 38020
rect 241336 6248 241388 6254
rect 241336 6190 241388 6196
rect 239588 4140 239640 4146
rect 239588 4082 239640 4088
rect 240048 4140 240100 4146
rect 240048 4082 240100 4088
rect 236092 604 236144 610
rect 236092 546 236144 552
rect 237196 604 237248 610
rect 237196 546 237248 552
rect 237564 604 237616 610
rect 237564 546 237616 552
rect 238392 604 238444 610
rect 238392 546 238444 552
rect 237208 480 237236 546
rect 238404 480 238432 546
rect 239600 480 239628 4082
rect 241440 3330 241468 38014
rect 241532 8838 241560 43302
rect 243464 40118 243492 43316
rect 244568 40118 244596 43316
rect 245488 40934 245516 43316
rect 245672 43302 246422 43330
rect 247052 43302 247526 43330
rect 245476 40928 245528 40934
rect 245476 40870 245528 40876
rect 243452 40112 243504 40118
rect 243452 40054 243504 40060
rect 244188 40112 244240 40118
rect 244188 40054 244240 40060
rect 244556 40112 244608 40118
rect 244556 40054 244608 40060
rect 245476 40112 245528 40118
rect 245476 40054 245528 40060
rect 242164 27056 242216 27062
rect 242164 26998 242216 27004
rect 241520 8832 241572 8838
rect 241520 8774 241572 8780
rect 241980 5160 242032 5166
rect 241980 5102 242032 5108
rect 240784 3324 240836 3330
rect 240784 3266 240836 3272
rect 241428 3324 241480 3330
rect 241428 3266 241480 3272
rect 240796 480 240824 3266
rect 241992 480 242020 5102
rect 242176 3874 242204 26998
rect 243176 9580 243228 9586
rect 243176 9522 243228 9528
rect 242164 3868 242216 3874
rect 242164 3810 242216 3816
rect 243188 480 243216 9522
rect 244200 6118 244228 40054
rect 245488 9586 245516 40054
rect 245568 38140 245620 38146
rect 245568 38082 245620 38088
rect 245476 9580 245528 9586
rect 245476 9522 245528 9528
rect 244188 6112 244240 6118
rect 244188 6054 244240 6060
rect 244372 3732 244424 3738
rect 244372 3674 244424 3680
rect 244384 480 244412 3674
rect 245580 480 245608 38082
rect 245672 6662 245700 43302
rect 245752 26988 245804 26994
rect 245752 26930 245804 26936
rect 245660 6656 245712 6662
rect 245660 6598 245712 6604
rect 245764 3346 245792 26930
rect 247052 12102 247080 43302
rect 248432 42770 248460 43316
rect 248420 42764 248472 42770
rect 248420 42706 248472 42712
rect 249352 40186 249380 43316
rect 250470 43302 251128 43330
rect 249340 40180 249392 40186
rect 249340 40122 249392 40128
rect 248420 22976 248472 22982
rect 248420 22918 248472 22924
rect 247132 16108 247184 16114
rect 247132 16050 247184 16056
rect 247040 12096 247092 12102
rect 247040 12038 247092 12044
rect 247144 3346 247172 16050
rect 248432 3482 248460 22918
rect 250352 9648 250404 9654
rect 250352 9590 250404 9596
rect 248432 3454 249196 3482
rect 245764 3318 246804 3346
rect 247144 3318 248000 3346
rect 246776 480 246804 3318
rect 247972 480 248000 3318
rect 249168 480 249196 3454
rect 250364 480 250392 9590
rect 251100 6730 251128 43302
rect 251192 43302 251390 43330
rect 251192 8906 251220 43302
rect 252480 11898 252508 43316
rect 253414 43302 253888 43330
rect 252560 35352 252612 35358
rect 252560 35294 252612 35300
rect 252468 11892 252520 11898
rect 252468 11834 252520 11840
rect 251180 8900 251232 8906
rect 251180 8842 251232 8848
rect 251088 6724 251140 6730
rect 251088 6666 251140 6672
rect 251456 3732 251508 3738
rect 251456 3674 251508 3680
rect 251468 480 251496 3674
rect 252572 3398 252600 35294
rect 253860 21554 253888 43302
rect 254320 40118 254348 43316
rect 255424 42022 255452 43316
rect 256358 43302 256648 43330
rect 255412 42016 255464 42022
rect 255412 41958 255464 41964
rect 255964 40180 256016 40186
rect 255964 40122 256016 40128
rect 254308 40112 254360 40118
rect 254308 40054 254360 40060
rect 255228 40112 255280 40118
rect 255228 40054 255280 40060
rect 252652 21548 252704 21554
rect 252652 21490 252704 21496
rect 253848 21548 253900 21554
rect 253848 21490 253900 21496
rect 252560 3392 252612 3398
rect 252560 3334 252612 3340
rect 252664 480 252692 21490
rect 255044 4140 255096 4146
rect 255044 4082 255096 4088
rect 253848 3392 253900 3398
rect 253848 3334 253900 3340
rect 253860 480 253888 3334
rect 255056 480 255084 4082
rect 255240 3806 255268 40054
rect 255976 3874 256004 40122
rect 256516 13252 256568 13258
rect 256516 13194 256568 13200
rect 255964 3868 256016 3874
rect 255964 3810 256016 3816
rect 255228 3800 255280 3806
rect 255228 3742 255280 3748
rect 256528 3482 256556 13194
rect 256620 8974 256648 43302
rect 257264 41274 257292 43316
rect 258368 41954 258396 43316
rect 260852 43302 261326 43330
rect 258356 41948 258408 41954
rect 258356 41890 258408 41896
rect 257252 41268 257304 41274
rect 257252 41210 257304 41216
rect 257436 9648 257488 9654
rect 257436 9590 257488 9596
rect 256608 8968 256660 8974
rect 256608 8910 256660 8916
rect 256252 3454 256556 3482
rect 256252 480 256280 3454
rect 257448 480 257476 9590
rect 260852 5098 260880 43302
rect 262128 41948 262180 41954
rect 262128 41890 262180 41896
rect 260840 5092 260892 5098
rect 260840 5034 260892 5040
rect 262140 3398 262168 41890
rect 264256 39982 264284 43316
rect 265176 39982 265204 43316
rect 266188 43302 266294 43330
rect 267214 43302 267688 43330
rect 268318 43302 268976 43330
rect 264244 39976 264296 39982
rect 264244 39918 264296 39924
rect 265164 39976 265216 39982
rect 265164 39918 265216 39924
rect 263508 39432 263560 39438
rect 263508 39374 263560 39380
rect 263416 35352 263468 35358
rect 263416 35294 263468 35300
rect 261024 3392 261076 3398
rect 261024 3334 261076 3340
rect 262128 3392 262180 3398
rect 262128 3334 262180 3340
rect 262220 3392 262272 3398
rect 262220 3334 262272 3340
rect 259828 3324 259880 3330
rect 259828 3266 259880 3272
rect 258632 3188 258684 3194
rect 258632 3130 258684 3136
rect 258644 480 258672 3130
rect 259840 480 259868 3266
rect 261036 480 261064 3334
rect 262232 480 262260 3334
rect 263428 480 263456 35294
rect 263520 3398 263548 39374
rect 264980 28484 265032 28490
rect 264980 28426 265032 28432
rect 264612 8900 264664 8906
rect 264612 8842 264664 8848
rect 263508 3392 263560 3398
rect 263508 3334 263560 3340
rect 264624 480 264652 8842
rect 264992 3482 265020 28426
rect 266188 6662 266216 43302
rect 266176 6656 266228 6662
rect 266176 6598 266228 6604
rect 267004 6044 267056 6050
rect 267004 5986 267056 5992
rect 264992 3454 265848 3482
rect 265820 480 265848 3454
rect 267016 480 267044 5986
rect 267660 5098 267688 43302
rect 268948 29646 268976 43302
rect 269224 40118 269252 43316
rect 270144 41342 270172 43316
rect 271262 43302 271828 43330
rect 274206 43302 274588 43330
rect 270132 41336 270184 41342
rect 270132 41278 270184 41284
rect 269212 40112 269264 40118
rect 269212 40054 269264 40060
rect 270408 40112 270460 40118
rect 270408 40054 270460 40060
rect 269028 32496 269080 32502
rect 269028 32438 269080 32444
rect 268936 29640 268988 29646
rect 268936 29582 268988 29588
rect 267648 5092 267700 5098
rect 267648 5034 267700 5040
rect 269040 3262 269068 32438
rect 269120 17536 269172 17542
rect 269120 17478 269172 17484
rect 269132 3482 269160 17478
rect 270420 16114 270448 40054
rect 270500 32564 270552 32570
rect 270500 32506 270552 32512
rect 270408 16108 270460 16114
rect 270408 16050 270460 16056
rect 269132 3454 269344 3482
rect 268108 3256 268160 3262
rect 268108 3198 268160 3204
rect 269028 3256 269080 3262
rect 269028 3198 269080 3204
rect 268120 480 268148 3198
rect 269316 480 269344 3454
rect 270512 480 270540 32506
rect 271800 31142 271828 43302
rect 271788 31136 271840 31142
rect 271788 31078 271840 31084
rect 274560 6594 274588 43302
rect 276032 43302 276230 43330
rect 278070 43302 278728 43330
rect 276032 29714 276060 43302
rect 276020 29708 276072 29714
rect 276020 29650 276072 29656
rect 275284 9444 275336 9450
rect 275284 9386 275336 9392
rect 272892 6588 272944 6594
rect 272892 6530 272944 6536
rect 274548 6588 274600 6594
rect 274548 6530 274600 6536
rect 271696 5092 271748 5098
rect 271696 5034 271748 5040
rect 271708 480 271736 5034
rect 272904 480 272932 6530
rect 274088 5024 274140 5030
rect 274088 4966 274140 4972
rect 274100 480 274128 4966
rect 275296 480 275324 9386
rect 277676 5976 277728 5982
rect 277676 5918 277728 5924
rect 276480 3256 276532 3262
rect 276480 3198 276532 3204
rect 276492 480 276520 3198
rect 277688 480 277716 5918
rect 278700 5030 278728 43302
rect 279160 40118 279188 43316
rect 279424 41472 279476 41478
rect 279424 41414 279476 41420
rect 279148 40112 279200 40118
rect 279148 40054 279200 40060
rect 278872 9308 278924 9314
rect 278872 9250 278924 9256
rect 278688 5024 278740 5030
rect 278688 4966 278740 4972
rect 278884 480 278912 9250
rect 279436 4078 279464 41414
rect 280068 40112 280120 40118
rect 280068 40054 280120 40060
rect 280080 31346 280108 40054
rect 280068 31340 280120 31346
rect 280068 31282 280120 31288
rect 280160 24200 280212 24206
rect 280160 24142 280212 24148
rect 279976 6520 280028 6526
rect 279976 6462 280028 6468
rect 279424 4072 279476 4078
rect 279424 4014 279476 4020
rect 279988 2666 280016 6462
rect 280066 4040 280122 4049
rect 280066 3975 280122 3984
rect 280080 2854 280108 3975
rect 280068 2848 280120 2854
rect 280068 2790 280120 2796
rect 279988 2638 280108 2666
rect 280080 480 280108 2638
rect 280172 610 280200 24142
rect 280632 20058 280660 43438
rect 281000 38010 281028 43316
rect 281092 38078 281120 59599
rect 281080 38072 281132 38078
rect 281080 38014 281132 38020
rect 280988 38004 281040 38010
rect 280988 37946 281040 37952
rect 280896 36508 280948 36514
rect 280896 36450 280948 36456
rect 280908 32502 280936 36450
rect 280896 32496 280948 32502
rect 280896 32438 280948 32444
rect 281184 25702 281212 84351
rect 281172 25696 281224 25702
rect 281172 25638 281224 25644
rect 280620 20052 280672 20058
rect 280620 19994 280672 20000
rect 281276 14618 281304 138479
rect 281368 135425 281396 154527
rect 281354 135416 281410 135425
rect 281354 135351 281410 135360
rect 281356 125520 281408 125526
rect 281356 125462 281408 125468
rect 281368 112402 281396 125462
rect 281552 124953 281580 461586
rect 281632 394732 281684 394738
rect 281632 394674 281684 394680
rect 281644 129305 281672 394674
rect 281908 336796 281960 336802
rect 281908 336738 281960 336744
rect 281816 268456 281868 268462
rect 281816 268398 281868 268404
rect 281724 266960 281776 266966
rect 281724 266902 281776 266908
rect 281630 129296 281686 129305
rect 281630 129231 281686 129240
rect 281538 124944 281594 124953
rect 281538 124879 281594 124888
rect 281356 112396 281408 112402
rect 281356 112338 281408 112344
rect 281356 106548 281408 106554
rect 281356 106490 281408 106496
rect 281368 94518 281396 106490
rect 281630 104952 281686 104961
rect 281630 104887 281686 104896
rect 281356 94512 281408 94518
rect 281356 94454 281408 94460
rect 281448 85060 281500 85066
rect 281448 85002 281500 85008
rect 281356 84924 281408 84930
rect 281356 84866 281408 84872
rect 281368 75342 281396 84866
rect 281356 75336 281408 75342
rect 281356 75278 281408 75284
rect 281460 75206 281488 85002
rect 281448 75200 281500 75206
rect 281448 75142 281500 75148
rect 281448 67448 281500 67454
rect 281448 67390 281500 67396
rect 281356 65476 281408 65482
rect 281356 65418 281408 65424
rect 281368 52766 281396 65418
rect 281356 52760 281408 52766
rect 281356 52702 281408 52708
rect 281460 51134 281488 67390
rect 281538 65376 281594 65385
rect 281538 65311 281594 65320
rect 281448 51128 281500 51134
rect 281448 51070 281500 51076
rect 281356 51060 281408 51066
rect 281356 51002 281408 51008
rect 281368 50946 281396 51002
rect 281368 50918 281488 50946
rect 281356 48272 281408 48278
rect 281356 48214 281408 48220
rect 281368 36514 281396 48214
rect 281460 36718 281488 50918
rect 281552 38146 281580 65311
rect 281540 38140 281592 38146
rect 281540 38082 281592 38088
rect 281448 36712 281500 36718
rect 281448 36654 281500 36660
rect 281540 36644 281592 36650
rect 281540 36586 281592 36592
rect 281356 36508 281408 36514
rect 281356 36450 281408 36456
rect 281264 14612 281316 14618
rect 281264 14554 281316 14560
rect 281552 4214 281580 36586
rect 281644 18834 281672 104887
rect 281632 18828 281684 18834
rect 281632 18770 281684 18776
rect 281540 4208 281592 4214
rect 281540 4150 281592 4156
rect 281540 4072 281592 4078
rect 281540 4014 281592 4020
rect 281552 3262 281580 4014
rect 281736 3942 281764 266902
rect 281828 6798 281856 268398
rect 281920 83609 281948 336738
rect 282276 267164 282328 267170
rect 282276 267106 282328 267112
rect 282000 266824 282052 266830
rect 282000 266766 282052 266772
rect 282012 258738 282040 266766
rect 282184 263492 282236 263498
rect 282184 263434 282236 263440
rect 282000 258732 282052 258738
rect 282000 258674 282052 258680
rect 282196 238066 282224 263434
rect 282288 257378 282316 267106
rect 282460 266756 282512 266762
rect 282460 266698 282512 266704
rect 282368 266620 282420 266626
rect 282368 266562 282420 266568
rect 282380 261662 282408 266562
rect 282472 263498 282500 266698
rect 282460 263492 282512 263498
rect 282460 263434 282512 263440
rect 282368 261656 282420 261662
rect 282368 261598 282420 261604
rect 282276 257372 282328 257378
rect 282276 257314 282328 257320
rect 282184 238060 282236 238066
rect 282184 238002 282236 238008
rect 282932 237402 282960 692786
rect 282840 237374 282960 237402
rect 281998 185872 282054 185881
rect 281998 185807 282054 185816
rect 281906 83600 281962 83609
rect 281906 83535 281962 83544
rect 281906 62928 281962 62937
rect 281906 62863 281962 62872
rect 281920 11966 281948 62863
rect 282012 39438 282040 185807
rect 282184 127628 282236 127634
rect 282184 127570 282236 127576
rect 282090 76256 282146 76265
rect 282090 76191 282146 76200
rect 282000 39432 282052 39438
rect 282000 39374 282052 39380
rect 282104 25770 282132 76191
rect 282092 25764 282144 25770
rect 282092 25706 282144 25712
rect 281908 11960 281960 11966
rect 281908 11902 281960 11908
rect 281816 6792 281868 6798
rect 281816 6734 281868 6740
rect 282196 4078 282224 127570
rect 282366 92304 282422 92313
rect 282366 92239 282422 92248
rect 282274 51232 282330 51241
rect 282274 51167 282330 51176
rect 282288 21486 282316 51167
rect 282380 33930 282408 92239
rect 282840 52465 282868 237374
rect 282918 235648 282974 235657
rect 282918 235583 282974 235592
rect 282826 52456 282882 52465
rect 282826 52391 282882 52400
rect 282368 33924 282420 33930
rect 282368 33866 282420 33872
rect 282276 21480 282328 21486
rect 282276 21422 282328 21428
rect 282932 7954 282960 235583
rect 283024 209681 283052 700538
rect 283852 692850 283880 703520
rect 287704 700528 287756 700534
rect 287704 700470 287756 700476
rect 283840 692844 283892 692850
rect 283840 692786 283892 692792
rect 284944 626612 284996 626618
rect 284944 626554 284996 626560
rect 283380 278044 283432 278050
rect 283380 277986 283432 277992
rect 283288 268184 283340 268190
rect 283288 268126 283340 268132
rect 283104 266688 283156 266694
rect 283104 266630 283156 266636
rect 283116 258806 283144 266630
rect 283194 261760 283250 261769
rect 283194 261695 283250 261704
rect 283208 260914 283236 261695
rect 283196 260908 283248 260914
rect 283196 260850 283248 260856
rect 283104 258800 283156 258806
rect 283104 258742 283156 258748
rect 283102 253056 283158 253065
rect 283102 252991 283158 253000
rect 283010 209672 283066 209681
rect 283010 209607 283066 209616
rect 283010 193216 283066 193225
rect 283010 193151 283066 193160
rect 283024 24478 283052 193151
rect 283116 43722 283144 252991
rect 283194 241360 283250 241369
rect 283194 241295 283250 241304
rect 283208 52601 283236 241295
rect 283300 179897 283328 268126
rect 283286 179888 283342 179897
rect 283286 179823 283342 179832
rect 283392 161242 283420 277986
rect 283472 273964 283524 273970
rect 283472 273906 283524 273912
rect 283484 191593 283512 273906
rect 284392 267776 284444 267782
rect 284392 267718 284444 267724
rect 283564 266552 283616 266558
rect 283564 266494 283616 266500
rect 283576 256018 283604 266494
rect 284300 265804 284352 265810
rect 284300 265746 284352 265752
rect 283564 256012 283616 256018
rect 283564 255954 283616 255960
rect 284114 251696 284170 251705
rect 284114 251631 284170 251640
rect 284128 251258 284156 251631
rect 284116 251252 284168 251258
rect 284116 251194 284168 251200
rect 284208 251184 284260 251190
rect 284208 251126 284260 251132
rect 284220 250073 284248 251126
rect 284206 250064 284262 250073
rect 284206 249999 284262 250008
rect 284206 248704 284262 248713
rect 284206 248639 284262 248648
rect 284220 248470 284248 248639
rect 284208 248464 284260 248470
rect 284208 248406 284260 248412
rect 284206 245712 284262 245721
rect 284206 245647 284208 245656
rect 284260 245647 284262 245656
rect 284208 245618 284260 245624
rect 284206 244352 284262 244361
rect 284206 244287 284208 244296
rect 284260 244287 284262 244296
rect 284208 244258 284260 244264
rect 283562 241496 283618 241505
rect 283562 241431 283618 241440
rect 283576 231985 283604 241431
rect 283840 238740 283892 238746
rect 283840 238682 283892 238688
rect 283852 238377 283880 238682
rect 283838 238368 283894 238377
rect 283838 238303 283894 238312
rect 283838 234832 283894 234841
rect 283838 234767 283894 234776
rect 283852 232121 283880 234767
rect 284206 234016 284262 234025
rect 284206 233951 284262 233960
rect 284220 233306 284248 233951
rect 284208 233300 284260 233306
rect 284208 233242 284260 233248
rect 283838 232112 283894 232121
rect 283838 232047 283894 232056
rect 283562 231976 283618 231985
rect 283562 231911 283618 231920
rect 284116 228608 284168 228614
rect 284116 228550 284168 228556
rect 284128 228313 284156 228550
rect 284114 228304 284170 228313
rect 284114 228239 284170 228248
rect 284206 226672 284262 226681
rect 284206 226607 284262 226616
rect 284220 226370 284248 226607
rect 284208 226364 284260 226370
rect 284208 226306 284260 226312
rect 284206 225312 284262 225321
rect 284206 225247 284262 225256
rect 284220 225010 284248 225247
rect 284208 225004 284260 225010
rect 284208 224946 284260 224952
rect 284206 217968 284262 217977
rect 284206 217903 284262 217912
rect 284220 216714 284248 217903
rect 284208 216708 284260 216714
rect 284208 216650 284260 216656
rect 284206 216608 284262 216617
rect 284206 216543 284262 216552
rect 284220 215354 284248 216543
rect 284208 215348 284260 215354
rect 284208 215290 284260 215296
rect 284206 213616 284262 213625
rect 284206 213551 284262 213560
rect 284220 212566 284248 213551
rect 284208 212560 284260 212566
rect 284208 212502 284260 212508
rect 284206 212256 284262 212265
rect 284206 212191 284262 212200
rect 284220 211206 284248 212191
rect 284208 211200 284260 211206
rect 284208 211142 284260 211148
rect 284114 207904 284170 207913
rect 284114 207839 284170 207848
rect 284128 207058 284156 207839
rect 284116 207052 284168 207058
rect 284116 206994 284168 207000
rect 284206 204912 284262 204921
rect 284206 204847 284262 204856
rect 284220 204406 284248 204847
rect 284208 204400 284260 204406
rect 284208 204342 284260 204348
rect 284206 201920 284262 201929
rect 284206 201855 284262 201864
rect 284220 201550 284248 201855
rect 284208 201544 284260 201550
rect 284208 201486 284260 201492
rect 284206 198928 284262 198937
rect 284206 198863 284262 198872
rect 284220 198762 284248 198863
rect 284208 198756 284260 198762
rect 284208 198698 284260 198704
rect 283562 197568 283618 197577
rect 283562 197503 283618 197512
rect 283470 191584 283526 191593
rect 283470 191519 283526 191528
rect 283300 161214 283420 161242
rect 283300 156505 283328 161214
rect 283378 161120 283434 161129
rect 283378 161055 283434 161064
rect 283392 160138 283420 161055
rect 283380 160132 283432 160138
rect 283380 160074 283432 160080
rect 283286 156496 283342 156505
rect 283286 156431 283342 156440
rect 283378 152144 283434 152153
rect 283378 152079 283434 152088
rect 283392 126993 283420 152079
rect 283576 127634 283604 197503
rect 284206 194576 284262 194585
rect 284206 194511 284262 194520
rect 284220 193254 284248 194511
rect 284208 193248 284260 193254
rect 284208 193190 284260 193196
rect 283838 192536 283894 192545
rect 283838 192471 283894 192480
rect 283852 180441 283880 192471
rect 284206 188864 284262 188873
rect 284206 188799 284262 188808
rect 284220 187746 284248 188799
rect 284208 187740 284260 187746
rect 284208 187682 284260 187688
rect 283930 184512 283986 184521
rect 283930 184447 283986 184456
rect 283838 180432 283894 180441
rect 283838 180367 283894 180376
rect 283838 165472 283894 165481
rect 283838 165407 283894 165416
rect 283852 164286 283880 165407
rect 283840 164280 283892 164286
rect 283840 164222 283892 164228
rect 283838 163840 283894 163849
rect 283838 163775 283894 163784
rect 283852 162926 283880 163775
rect 283840 162920 283892 162926
rect 283840 162862 283892 162868
rect 283840 150408 283892 150414
rect 283840 150350 283892 150356
rect 283852 149433 283880 150350
rect 283838 149424 283894 149433
rect 283838 149359 283894 149368
rect 283840 144900 283892 144906
rect 283840 144842 283892 144848
rect 283852 144809 283880 144842
rect 283838 144800 283894 144809
rect 283838 144735 283894 144744
rect 283838 143440 283894 143449
rect 283838 143375 283894 143384
rect 283852 142186 283880 143375
rect 283840 142180 283892 142186
rect 283840 142122 283892 142128
rect 283746 137728 283802 137737
rect 283746 137663 283802 137672
rect 283760 136678 283788 137663
rect 283748 136672 283800 136678
rect 283748 136614 283800 136620
rect 283564 127628 283616 127634
rect 283564 127570 283616 127576
rect 283470 127392 283526 127401
rect 283470 127327 283526 127336
rect 283378 126984 283434 126993
rect 283378 126919 283434 126928
rect 283378 126032 283434 126041
rect 283378 125967 283434 125976
rect 283286 52864 283342 52873
rect 283286 52799 283342 52808
rect 283194 52592 283250 52601
rect 283194 52527 283250 52536
rect 283300 49178 283328 52799
rect 283208 49150 283328 49178
rect 283104 43716 283156 43722
rect 283104 43658 283156 43664
rect 283208 38214 283236 49150
rect 283196 38208 283248 38214
rect 283196 38150 283248 38156
rect 283012 24472 283064 24478
rect 283012 24414 283064 24420
rect 283392 13258 283420 125967
rect 283484 23050 283512 127327
rect 283838 121408 283894 121417
rect 283838 121343 283894 121352
rect 283852 120154 283880 121343
rect 283840 120148 283892 120154
rect 283840 120090 283892 120096
rect 283654 118688 283710 118697
rect 283654 118623 283710 118632
rect 283668 117366 283696 118623
rect 283656 117360 283708 117366
rect 283656 117302 283708 117308
rect 283562 117056 283618 117065
rect 283562 116991 283618 117000
rect 283472 23044 283524 23050
rect 283472 22986 283524 22992
rect 283576 16182 283604 116991
rect 283746 112704 283802 112713
rect 283746 112639 283802 112648
rect 283760 111858 283788 112639
rect 283748 111852 283800 111858
rect 283748 111794 283800 111800
rect 283838 104000 283894 104009
rect 283838 103935 283894 103944
rect 283852 103562 283880 103935
rect 283840 103556 283892 103562
rect 283840 103498 283892 103504
rect 283654 99648 283710 99657
rect 283654 99583 283710 99592
rect 283668 99414 283696 99583
rect 283656 99408 283708 99414
rect 283656 99350 283708 99356
rect 283840 98048 283892 98054
rect 283838 98016 283840 98025
rect 283892 98016 283894 98025
rect 283838 97951 283894 97960
rect 283746 96656 283802 96665
rect 283746 96591 283802 96600
rect 283654 81968 283710 81977
rect 283654 81903 283710 81912
rect 283668 81462 283696 81903
rect 283656 81456 283708 81462
rect 283656 81398 283708 81404
rect 283654 80608 283710 80617
rect 283654 80543 283710 80552
rect 283564 16176 283616 16182
rect 283564 16118 283616 16124
rect 283380 13252 283432 13258
rect 283380 13194 283432 13200
rect 283012 12028 283064 12034
rect 283012 11970 283064 11976
rect 282920 7948 282972 7954
rect 282920 7890 282972 7896
rect 282460 4208 282512 4214
rect 282460 4150 282512 4156
rect 282184 4072 282236 4078
rect 282184 4014 282236 4020
rect 281724 3936 281776 3942
rect 281724 3878 281776 3884
rect 281540 3256 281592 3262
rect 281540 3198 281592 3204
rect 280160 604 280212 610
rect 280160 546 280212 552
rect 281264 604 281316 610
rect 281264 546 281316 552
rect 281276 480 281304 546
rect 282472 480 282500 4150
rect 283024 3380 283052 11970
rect 283668 5166 283696 80543
rect 283760 35358 283788 96591
rect 283838 95296 283894 95305
rect 283838 95231 283840 95240
rect 283892 95231 283894 95240
rect 283840 95202 283892 95208
rect 283840 93832 283892 93838
rect 283840 93774 283892 93780
rect 283852 93673 283880 93774
rect 283838 93664 283894 93673
rect 283838 93599 283894 93608
rect 283840 89684 283892 89690
rect 283840 89626 283892 89632
rect 283852 89321 283880 89626
rect 283838 89312 283894 89321
rect 283838 89247 283894 89256
rect 283838 87952 283894 87961
rect 283838 87887 283894 87896
rect 283852 87038 283880 87887
rect 283840 87032 283892 87038
rect 283840 86974 283892 86980
rect 283838 86320 283894 86329
rect 283838 86255 283894 86264
rect 283852 85610 283880 86255
rect 283840 85604 283892 85610
rect 283840 85546 283892 85552
rect 283838 68912 283894 68921
rect 283838 68847 283894 68856
rect 283852 67658 283880 68847
rect 283840 67652 283892 67658
rect 283840 67594 283892 67600
rect 283838 64560 283894 64569
rect 283838 64495 283894 64504
rect 283852 63578 283880 64495
rect 283840 63572 283892 63578
rect 283840 63514 283892 63520
rect 283840 62076 283892 62082
rect 283840 62018 283892 62024
rect 283852 61577 283880 62018
rect 283838 61568 283894 61577
rect 283838 61503 283894 61512
rect 283838 58576 283894 58585
rect 283838 58511 283894 58520
rect 283852 58002 283880 58511
rect 283840 57996 283892 58002
rect 283840 57938 283892 57944
rect 283838 46880 283894 46889
rect 283838 46815 283894 46824
rect 283852 45626 283880 46815
rect 283840 45620 283892 45626
rect 283840 45562 283892 45568
rect 283838 45520 283894 45529
rect 283838 45455 283894 45464
rect 283852 44198 283880 45455
rect 283840 44192 283892 44198
rect 283840 44134 283892 44140
rect 283748 35352 283800 35358
rect 283748 35294 283800 35300
rect 283944 27062 283972 184447
rect 284206 182880 284262 182889
rect 284206 182815 284262 182824
rect 284220 182238 284248 182815
rect 284208 182232 284260 182238
rect 284208 182174 284260 182180
rect 284206 177168 284262 177177
rect 284206 177103 284262 177112
rect 284220 176730 284248 177103
rect 284208 176724 284260 176730
rect 284208 176666 284260 176672
rect 284206 174176 284262 174185
rect 284206 174111 284262 174120
rect 284220 173942 284248 174111
rect 284208 173936 284260 173942
rect 284208 173878 284260 173884
rect 284206 171184 284262 171193
rect 284206 171119 284208 171128
rect 284260 171119 284262 171128
rect 284208 171090 284260 171096
rect 284022 153776 284078 153785
rect 284022 153711 284078 153720
rect 284036 153270 284064 153711
rect 284024 153264 284076 153270
rect 284024 153206 284076 153212
rect 284208 142112 284260 142118
rect 284206 142080 284208 142089
rect 284260 142080 284262 142089
rect 284206 142015 284262 142024
rect 284206 136096 284262 136105
rect 284206 136031 284262 136040
rect 284220 135318 284248 136031
rect 284208 135312 284260 135318
rect 284208 135254 284260 135260
rect 284022 109712 284078 109721
rect 284022 109647 284078 109656
rect 284036 109070 284064 109647
rect 284024 109064 284076 109070
rect 284024 109006 284076 109012
rect 284022 108352 284078 108361
rect 284022 108287 284078 108296
rect 284036 107710 284064 108287
rect 284024 107704 284076 107710
rect 284024 107646 284076 107652
rect 284022 106992 284078 107001
rect 284022 106927 284078 106936
rect 284036 106350 284064 106927
rect 284024 106344 284076 106350
rect 284024 106286 284076 106292
rect 284206 101008 284262 101017
rect 284206 100943 284262 100952
rect 284220 100774 284248 100943
rect 284208 100768 284260 100774
rect 284208 100710 284260 100716
rect 284022 90944 284078 90953
rect 284022 90879 284078 90888
rect 284036 89758 284064 90879
rect 284024 89752 284076 89758
rect 284024 89694 284076 89700
rect 284206 78976 284262 78985
rect 284206 78911 284262 78920
rect 284220 78742 284248 78911
rect 284208 78736 284260 78742
rect 284208 78678 284260 78684
rect 284206 74624 284262 74633
rect 284206 74559 284208 74568
rect 284260 74559 284262 74568
rect 284208 74530 284260 74536
rect 284206 71904 284262 71913
rect 284206 71839 284262 71848
rect 284220 71806 284248 71839
rect 284208 71800 284260 71806
rect 284208 71742 284260 71748
rect 283932 27056 283984 27062
rect 283932 26998 283984 27004
rect 283656 5160 283708 5166
rect 283656 5102 283708 5108
rect 284312 3482 284340 265746
rect 284404 6050 284432 267718
rect 284576 265396 284628 265402
rect 284576 265338 284628 265344
rect 284484 264512 284536 264518
rect 284484 264454 284536 264460
rect 284392 6044 284444 6050
rect 284392 5986 284444 5992
rect 284496 3738 284524 264454
rect 284588 6866 284616 265338
rect 284668 264580 284720 264586
rect 284668 264522 284720 264528
rect 284680 41478 284708 264522
rect 284668 41472 284720 41478
rect 284668 41414 284720 41420
rect 284956 39778 284984 626554
rect 285036 509312 285088 509318
rect 285036 509254 285088 509260
rect 285048 41993 285076 509254
rect 286324 404388 286376 404394
rect 286324 404330 286376 404336
rect 285128 345092 285180 345098
rect 285128 345034 285180 345040
rect 285140 42702 285168 345034
rect 285956 269884 286008 269890
rect 285956 269826 286008 269832
rect 285680 269612 285732 269618
rect 285680 269554 285732 269560
rect 285218 263936 285274 263945
rect 285218 263871 285274 263880
rect 285128 42696 285180 42702
rect 285128 42638 285180 42644
rect 285034 41984 285090 41993
rect 285034 41919 285090 41928
rect 284944 39772 284996 39778
rect 284944 39714 284996 39720
rect 284576 6860 284628 6866
rect 284576 6802 284628 6808
rect 285232 3738 285260 263871
rect 285312 169788 285364 169794
rect 285312 169730 285364 169736
rect 285324 42022 285352 169730
rect 285312 42016 285364 42022
rect 285312 41958 285364 41964
rect 284484 3732 284536 3738
rect 284484 3674 284536 3680
rect 285220 3732 285272 3738
rect 285220 3674 285272 3680
rect 284312 3454 284800 3482
rect 283024 3352 283696 3380
rect 283668 480 283696 3352
rect 284772 480 284800 3454
rect 285692 3398 285720 269554
rect 285772 264648 285824 264654
rect 285772 264590 285824 264596
rect 285784 4010 285812 264590
rect 285864 263084 285916 263090
rect 285864 263026 285916 263032
rect 285772 4004 285824 4010
rect 285772 3946 285824 3952
rect 285680 3392 285732 3398
rect 285680 3334 285732 3340
rect 285876 3330 285904 263026
rect 285968 42226 285996 269826
rect 286048 269136 286100 269142
rect 286048 269078 286100 269084
rect 285956 42220 286008 42226
rect 285956 42162 286008 42168
rect 286060 42158 286088 269078
rect 286140 265532 286192 265538
rect 286140 265474 286192 265480
rect 286152 42430 286180 265474
rect 286232 100768 286284 100774
rect 286232 100710 286284 100716
rect 286140 42424 286192 42430
rect 286140 42366 286192 42372
rect 286244 42362 286272 100710
rect 286336 42906 286364 404330
rect 286416 392012 286468 392018
rect 286416 391954 286468 391960
rect 286324 42900 286376 42906
rect 286324 42842 286376 42848
rect 286428 42770 286456 391954
rect 286508 282192 286560 282198
rect 286508 282134 286560 282140
rect 286520 228614 286548 282134
rect 287152 269680 287204 269686
rect 287152 269622 287204 269628
rect 287060 264988 287112 264994
rect 287060 264930 287112 264936
rect 286600 262812 286652 262818
rect 286600 262754 286652 262760
rect 286612 252550 286640 262754
rect 286600 252544 286652 252550
rect 286600 252486 286652 252492
rect 286508 228608 286560 228614
rect 286508 228550 286560 228556
rect 286508 81456 286560 81462
rect 286508 81398 286560 81404
rect 286416 42764 286468 42770
rect 286416 42706 286468 42712
rect 286232 42356 286284 42362
rect 286232 42298 286284 42304
rect 286048 42152 286100 42158
rect 286048 42094 286100 42100
rect 285954 37904 286010 37913
rect 285954 37839 286010 37848
rect 285864 3324 285916 3330
rect 285864 3266 285916 3272
rect 285968 480 285996 37839
rect 286520 35902 286548 81398
rect 286508 35896 286560 35902
rect 286508 35838 286560 35844
rect 287072 3398 287100 264930
rect 287164 4146 287192 269622
rect 287244 269204 287296 269210
rect 287244 269146 287296 269152
rect 287256 42294 287284 269146
rect 287716 42498 287744 700470
rect 290464 700392 290516 700398
rect 290464 700334 290516 700340
rect 289820 269816 289872 269822
rect 289820 269758 289872 269764
rect 288532 269748 288584 269754
rect 288532 269690 288584 269696
rect 287888 267232 287940 267238
rect 287888 267174 287940 267180
rect 287796 266892 287848 266898
rect 287796 266834 287848 266840
rect 287808 44878 287836 266834
rect 287900 86290 287928 267174
rect 287978 266928 288034 266937
rect 287978 266863 288034 266872
rect 287992 243574 288020 266863
rect 288440 263560 288492 263566
rect 288440 263502 288492 263508
rect 287980 243568 288032 243574
rect 287980 243510 288032 243516
rect 287888 86284 287940 86290
rect 287888 86226 287940 86232
rect 287796 44872 287848 44878
rect 287796 44814 287848 44820
rect 287704 42492 287756 42498
rect 287704 42434 287756 42440
rect 287244 42288 287296 42294
rect 287244 42230 287296 42236
rect 287244 31340 287296 31346
rect 287244 31282 287296 31288
rect 287152 4140 287204 4146
rect 287152 4082 287204 4088
rect 287256 3482 287284 31282
rect 287164 3454 287284 3482
rect 288452 3482 288480 263502
rect 288544 5982 288572 269690
rect 288624 268388 288676 268394
rect 288624 268330 288676 268336
rect 288636 9654 288664 268330
rect 288716 266484 288768 266490
rect 288716 266426 288768 266432
rect 288728 41954 288756 266426
rect 288716 41948 288768 41954
rect 288716 41890 288768 41896
rect 288624 9648 288676 9654
rect 288624 9590 288676 9596
rect 289832 8906 289860 269758
rect 290476 93838 290504 700334
rect 300136 688634 300164 703520
rect 332520 700534 332548 703520
rect 332508 700528 332560 700534
rect 332508 700470 332560 700476
rect 348804 700466 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365116 703474
rect 348792 700460 348844 700466
rect 348792 700402 348844 700408
rect 319444 696992 319496 696998
rect 319444 696934 319496 696940
rect 299664 688628 299716 688634
rect 299664 688570 299716 688576
rect 300124 688628 300176 688634
rect 300124 688570 300176 688576
rect 299676 685930 299704 688570
rect 295984 685908 296036 685914
rect 295984 685850 296036 685856
rect 299584 685902 299704 685930
rect 293224 638988 293276 638994
rect 293224 638930 293276 638936
rect 291844 485852 291896 485858
rect 291844 485794 291896 485800
rect 290556 274712 290608 274718
rect 290556 274654 290608 274660
rect 290464 93832 290516 93838
rect 290464 93774 290516 93780
rect 289912 63572 289964 63578
rect 289912 63514 289964 63520
rect 289820 8900 289872 8906
rect 289820 8842 289872 8848
rect 288532 5976 288584 5982
rect 288532 5918 288584 5924
rect 288452 3454 289584 3482
rect 287060 3392 287112 3398
rect 287060 3334 287112 3340
rect 287164 480 287192 3454
rect 288348 3392 288400 3398
rect 288348 3334 288400 3340
rect 288360 480 288388 3334
rect 289556 480 289584 3454
rect 289924 3346 289952 63514
rect 290568 42634 290596 274654
rect 290556 42628 290608 42634
rect 290556 42570 290608 42576
rect 291856 39710 291884 485794
rect 291936 321632 291988 321638
rect 291936 321574 291988 321580
rect 291948 42566 291976 321574
rect 292580 182232 292632 182238
rect 292580 182174 292632 182180
rect 291936 42560 291988 42566
rect 291936 42502 291988 42508
rect 291844 39704 291896 39710
rect 291844 39646 291896 39652
rect 291200 16108 291252 16114
rect 291200 16050 291252 16056
rect 291212 3346 291240 16050
rect 292592 3346 292620 182174
rect 293236 42401 293264 638930
rect 294604 498228 294656 498234
rect 294604 498170 294656 498176
rect 293316 268524 293368 268530
rect 293316 268466 293368 268472
rect 293328 182170 293356 268466
rect 293316 182164 293368 182170
rect 293316 182106 293368 182112
rect 294616 42809 294644 498170
rect 294696 268592 294748 268598
rect 294696 268534 294748 268540
rect 294708 77246 294736 268534
rect 294696 77240 294748 77246
rect 294696 77182 294748 77188
rect 294602 42800 294658 42809
rect 294602 42735 294658 42744
rect 293222 42392 293278 42401
rect 293222 42327 293278 42336
rect 295996 39846 296024 685850
rect 299584 684486 299612 685902
rect 299572 684480 299624 684486
rect 299572 684422 299624 684428
rect 299940 666596 299992 666602
rect 299940 666538 299992 666544
rect 299952 659682 299980 666538
rect 299768 659654 299980 659682
rect 299768 647290 299796 659654
rect 313924 650072 313976 650078
rect 313924 650014 313976 650020
rect 299664 647284 299716 647290
rect 299664 647226 299716 647232
rect 299756 647284 299808 647290
rect 299756 647226 299808 647232
rect 299676 640422 299704 647226
rect 299664 640416 299716 640422
rect 299664 640358 299716 640364
rect 299756 640416 299808 640422
rect 299756 640358 299808 640364
rect 299768 630698 299796 640358
rect 299572 630692 299624 630698
rect 299572 630634 299624 630640
rect 299756 630692 299808 630698
rect 299756 630634 299808 630640
rect 299584 630578 299612 630634
rect 299584 630550 299704 630578
rect 299676 621058 299704 630550
rect 299676 621030 299796 621058
rect 299768 611386 299796 621030
rect 299572 611380 299624 611386
rect 299572 611322 299624 611328
rect 299756 611380 299808 611386
rect 299756 611322 299808 611328
rect 299584 611266 299612 611322
rect 299584 611238 299704 611266
rect 299676 608598 299704 611238
rect 299664 608592 299716 608598
rect 299664 608534 299716 608540
rect 299848 601724 299900 601730
rect 299848 601666 299900 601672
rect 299860 598942 299888 601666
rect 299848 598936 299900 598942
rect 299848 598878 299900 598884
rect 299940 589348 299992 589354
rect 299940 589290 299992 589296
rect 299952 582486 299980 589290
rect 299940 582480 299992 582486
rect 299940 582422 299992 582428
rect 299848 582344 299900 582350
rect 299848 582286 299900 582292
rect 299860 572642 299888 582286
rect 299676 572614 299888 572642
rect 299676 569945 299704 572614
rect 299662 569936 299718 569945
rect 299662 569871 299718 569880
rect 299570 560416 299626 560425
rect 299570 560351 299626 560360
rect 299584 553466 299612 560351
rect 299584 553438 299704 553466
rect 299676 550662 299704 553438
rect 299480 550656 299532 550662
rect 299480 550598 299532 550604
rect 299664 550656 299716 550662
rect 299664 550598 299716 550604
rect 299492 549273 299520 550598
rect 299294 549264 299350 549273
rect 299294 549199 299350 549208
rect 299478 549264 299534 549273
rect 299478 549199 299534 549208
rect 299308 543726 299336 549199
rect 299296 543720 299348 543726
rect 299296 543662 299348 543668
rect 299480 543720 299532 543726
rect 299480 543662 299532 543668
rect 299492 539594 299520 543662
rect 299492 539566 299612 539594
rect 299584 531350 299612 539566
rect 299572 531344 299624 531350
rect 299572 531286 299624 531292
rect 299756 531344 299808 531350
rect 299756 531286 299808 531292
rect 299768 524482 299796 531286
rect 299756 524476 299808 524482
rect 299756 524418 299808 524424
rect 299848 524408 299900 524414
rect 299848 524350 299900 524356
rect 299860 521665 299888 524350
rect 299662 521656 299718 521665
rect 299662 521591 299718 521600
rect 299846 521656 299902 521665
rect 299846 521591 299902 521600
rect 299676 512038 299704 521591
rect 299664 512032 299716 512038
rect 299664 511974 299716 511980
rect 299940 512032 299992 512038
rect 299940 511974 299992 511980
rect 299952 502382 299980 511974
rect 299756 502376 299808 502382
rect 299478 502344 299534 502353
rect 299478 502279 299534 502288
rect 299754 502344 299756 502353
rect 299940 502376 299992 502382
rect 299808 502344 299810 502353
rect 299940 502318 299992 502324
rect 299754 502279 299810 502288
rect 299492 492697 299520 502279
rect 299478 492688 299534 492697
rect 299478 492623 299534 492632
rect 299662 492688 299718 492697
rect 299662 492623 299664 492632
rect 299716 492623 299718 492632
rect 299664 492594 299716 492600
rect 299664 485784 299716 485790
rect 299664 485726 299716 485732
rect 299676 483018 299704 485726
rect 299676 482990 299796 483018
rect 299768 476134 299796 482990
rect 299572 476128 299624 476134
rect 299756 476128 299808 476134
rect 299624 476076 299704 476082
rect 299572 476070 299704 476076
rect 299756 476070 299808 476076
rect 299584 476054 299704 476070
rect 299676 473346 299704 476054
rect 299664 473340 299716 473346
rect 299664 473282 299716 473288
rect 299664 466404 299716 466410
rect 299664 466346 299716 466352
rect 299676 463706 299704 466346
rect 299676 463678 299796 463706
rect 299768 460902 299796 463678
rect 299388 460896 299440 460902
rect 299388 460838 299440 460844
rect 299756 460896 299808 460902
rect 299756 460838 299808 460844
rect 299400 451330 299428 460838
rect 299400 451302 299520 451330
rect 299492 449886 299520 451302
rect 299480 449880 299532 449886
rect 299480 449822 299532 449828
rect 299572 440292 299624 440298
rect 299572 440234 299624 440240
rect 299584 436830 299612 440234
rect 299572 436824 299624 436830
rect 299572 436766 299624 436772
rect 299572 423700 299624 423706
rect 299572 423642 299624 423648
rect 299584 422278 299612 423642
rect 299572 422272 299624 422278
rect 299572 422214 299624 422220
rect 299756 422272 299808 422278
rect 299756 422214 299808 422220
rect 299768 412729 299796 422214
rect 299478 412720 299534 412729
rect 299478 412655 299534 412664
rect 299754 412720 299810 412729
rect 299754 412655 299810 412664
rect 299492 412622 299520 412655
rect 299480 412616 299532 412622
rect 299480 412558 299532 412564
rect 299572 412616 299624 412622
rect 299572 412558 299624 412564
rect 299584 401606 299612 412558
rect 299204 401600 299256 401606
rect 299204 401542 299256 401548
rect 299572 401600 299624 401606
rect 299572 401542 299624 401548
rect 299216 392057 299244 401542
rect 299202 392048 299258 392057
rect 299202 391983 299258 391992
rect 299386 392048 299442 392057
rect 299386 391983 299442 391992
rect 299400 391950 299428 391983
rect 299388 391944 299440 391950
rect 299388 391886 299440 391892
rect 299572 389088 299624 389094
rect 299572 389030 299624 389036
rect 299584 379506 299612 389030
rect 299572 379500 299624 379506
rect 299572 379442 299624 379448
rect 299756 379500 299808 379506
rect 299756 379442 299808 379448
rect 299768 371906 299796 379442
rect 299768 371878 299888 371906
rect 299860 357542 299888 371878
rect 299848 357536 299900 357542
rect 299848 357478 299900 357484
rect 304356 357468 304408 357474
rect 304356 357410 304408 357416
rect 299756 356176 299808 356182
rect 299808 356124 299888 356130
rect 299756 356118 299888 356124
rect 299768 356102 299888 356118
rect 299860 354686 299888 356102
rect 299848 354680 299900 354686
rect 299848 354622 299900 354628
rect 299940 336796 299992 336802
rect 299940 336738 299992 336744
rect 299952 331378 299980 336738
rect 299860 331350 299980 331378
rect 299860 327146 299888 331350
rect 299756 327140 299808 327146
rect 299756 327082 299808 327088
rect 299848 327140 299900 327146
rect 299848 327082 299900 327088
rect 299768 318850 299796 327082
rect 299664 318844 299716 318850
rect 299664 318786 299716 318792
rect 299756 318844 299808 318850
rect 299756 318786 299808 318792
rect 299676 311982 299704 318786
rect 299664 311976 299716 311982
rect 299664 311918 299716 311924
rect 299756 311976 299808 311982
rect 299756 311918 299808 311924
rect 299768 302258 299796 311918
rect 299572 302252 299624 302258
rect 299572 302194 299624 302200
rect 299756 302252 299808 302258
rect 299756 302194 299808 302200
rect 299584 302138 299612 302194
rect 299584 302110 299704 302138
rect 299676 299470 299704 302110
rect 299664 299464 299716 299470
rect 299664 299406 299716 299412
rect 299756 289876 299808 289882
rect 299756 289818 299808 289824
rect 299768 282826 299796 289818
rect 299676 282798 299796 282826
rect 299676 273329 299704 282798
rect 299662 273320 299718 273329
rect 299662 273255 299718 273264
rect 299662 270600 299718 270609
rect 299662 270535 299718 270544
rect 298100 265464 298152 265470
rect 298100 265406 298152 265412
rect 296720 264172 296772 264178
rect 296720 264114 296772 264120
rect 295984 39840 296036 39846
rect 295984 39782 296036 39788
rect 295340 31204 295392 31210
rect 295340 31146 295392 31152
rect 294328 9172 294380 9178
rect 294328 9114 294380 9120
rect 289924 3318 290780 3346
rect 291212 3318 291976 3346
rect 292592 3318 293172 3346
rect 290752 480 290780 3318
rect 291948 480 291976 3318
rect 293144 480 293172 3318
rect 294340 480 294368 9114
rect 295352 3346 295380 31146
rect 296732 3398 296760 264114
rect 296812 261656 296864 261662
rect 296812 261598 296864 261604
rect 296720 3392 296772 3398
rect 295352 3318 295564 3346
rect 296720 3334 296772 3340
rect 295536 480 295564 3318
rect 296824 1442 296852 261598
rect 298112 3482 298140 265406
rect 299676 260846 299704 270535
rect 300860 264376 300912 264382
rect 300860 264318 300912 264324
rect 299480 260840 299532 260846
rect 299480 260782 299532 260788
rect 299664 260840 299716 260846
rect 299664 260782 299716 260788
rect 299492 251297 299520 260782
rect 299478 251288 299534 251297
rect 299478 251223 299534 251232
rect 299754 251288 299810 251297
rect 299754 251223 299810 251232
rect 299768 244202 299796 251223
rect 299676 244174 299796 244202
rect 299676 241505 299704 244174
rect 299478 241496 299534 241505
rect 299478 241431 299534 241440
rect 299662 241496 299718 241505
rect 299662 241431 299718 241440
rect 299492 231878 299520 241431
rect 299480 231872 299532 231878
rect 299480 231814 299532 231820
rect 299756 231872 299808 231878
rect 299756 231814 299808 231820
rect 299768 224890 299796 231814
rect 299676 224862 299796 224890
rect 299676 222193 299704 224862
rect 299478 222184 299534 222193
rect 299478 222119 299534 222128
rect 299662 222184 299718 222193
rect 299662 222119 299718 222128
rect 299492 212634 299520 222119
rect 299480 212628 299532 212634
rect 299480 212570 299532 212576
rect 299756 212628 299808 212634
rect 299756 212570 299808 212576
rect 299768 205578 299796 212570
rect 299676 205550 299796 205578
rect 299676 202842 299704 205550
rect 299664 202836 299716 202842
rect 299664 202778 299716 202784
rect 299756 193316 299808 193322
rect 299756 193258 299808 193264
rect 299768 186266 299796 193258
rect 299676 186238 299796 186266
rect 299676 183569 299704 186238
rect 299478 183560 299534 183569
rect 299478 183495 299534 183504
rect 299662 183560 299718 183569
rect 299662 183495 299718 183504
rect 299492 174010 299520 183495
rect 299480 174004 299532 174010
rect 299480 173946 299532 173952
rect 299756 174004 299808 174010
rect 299756 173946 299808 173952
rect 299768 166954 299796 173946
rect 299676 166926 299796 166954
rect 299676 164218 299704 166926
rect 299480 164212 299532 164218
rect 299480 164154 299532 164160
rect 299664 164212 299716 164218
rect 299664 164154 299716 164160
rect 299492 154601 299520 164154
rect 299478 154592 299534 154601
rect 299478 154527 299534 154536
rect 299754 154592 299810 154601
rect 299754 154527 299810 154536
rect 299768 147642 299796 154527
rect 299676 147614 299796 147642
rect 299676 140026 299704 147614
rect 299492 139998 299704 140026
rect 299492 135289 299520 139998
rect 299478 135280 299534 135289
rect 299478 135215 299534 135224
rect 299754 135280 299810 135289
rect 299754 135215 299810 135224
rect 299768 128330 299796 135215
rect 299676 128302 299796 128330
rect 299676 120714 299704 128302
rect 299492 120686 299704 120714
rect 299492 115977 299520 120686
rect 299478 115968 299534 115977
rect 299478 115903 299534 115912
rect 299754 115968 299810 115977
rect 299754 115903 299810 115912
rect 299768 109018 299796 115903
rect 299676 108990 299796 109018
rect 299676 101454 299704 108990
rect 299664 101448 299716 101454
rect 299664 101390 299716 101396
rect 299664 99340 299716 99346
rect 299664 99282 299716 99288
rect 299676 96642 299704 99282
rect 299676 96614 299796 96642
rect 299768 89706 299796 96614
rect 299676 89678 299796 89706
rect 299676 86970 299704 89678
rect 299664 86964 299716 86970
rect 299664 86906 299716 86912
rect 299664 77308 299716 77314
rect 299664 77250 299716 77256
rect 299676 67590 299704 77250
rect 299664 67584 299716 67590
rect 299664 67526 299716 67532
rect 299664 60988 299716 60994
rect 299664 60930 299716 60936
rect 299676 51082 299704 60930
rect 299676 51054 299796 51082
rect 299768 39914 299796 51054
rect 299756 39908 299808 39914
rect 299756 39850 299808 39856
rect 299480 11824 299532 11830
rect 299480 11766 299532 11772
rect 299492 3482 299520 11766
rect 300872 3482 300900 264318
rect 304264 260908 304316 260914
rect 304264 260850 304316 260856
rect 302240 248464 302292 248470
rect 302240 248406 302292 248412
rect 302252 3482 302280 248406
rect 304276 16114 304304 260850
rect 304368 251190 304396 357410
rect 305000 267096 305052 267102
rect 305000 267038 305052 267044
rect 304356 251184 304408 251190
rect 304356 251126 304408 251132
rect 304356 204332 304408 204338
rect 304356 204274 304408 204280
rect 304368 62082 304396 204274
rect 304356 62076 304408 62082
rect 304356 62018 304408 62024
rect 304264 16108 304316 16114
rect 304264 16050 304316 16056
rect 303804 9580 303856 9586
rect 303804 9522 303856 9528
rect 298112 3454 299152 3482
rect 299492 3454 300348 3482
rect 300872 3454 301452 3482
rect 302252 3454 302648 3482
rect 297916 3392 297968 3398
rect 297916 3334 297968 3340
rect 296732 1414 296852 1442
rect 296732 480 296760 1414
rect 297928 480 297956 3334
rect 299124 480 299152 3454
rect 300320 480 300348 3454
rect 301424 480 301452 3454
rect 302620 480 302648 3454
rect 303816 480 303844 9522
rect 305012 480 305040 267038
rect 306380 258800 306432 258806
rect 306380 258742 306432 258748
rect 305644 204400 305696 204406
rect 305644 204342 305696 204348
rect 305656 50386 305684 204342
rect 305644 50380 305696 50386
rect 305644 50322 305696 50328
rect 306196 6112 306248 6118
rect 306196 6054 306248 6060
rect 306208 480 306236 6054
rect 306392 3482 306420 258742
rect 311900 245676 311952 245682
rect 311900 245618 311952 245624
rect 308404 233300 308456 233306
rect 308404 233242 308456 233248
rect 307760 31272 307812 31278
rect 307760 31214 307812 31220
rect 307772 3482 307800 31214
rect 308416 11830 308444 233242
rect 308496 133952 308548 133958
rect 308496 133894 308548 133900
rect 308508 89690 308536 133894
rect 308496 89684 308548 89690
rect 308496 89626 308548 89632
rect 310520 44872 310572 44878
rect 310520 44814 310572 44820
rect 309140 16040 309192 16046
rect 309140 15982 309192 15988
rect 308404 11824 308456 11830
rect 308404 11766 308456 11772
rect 309152 3482 309180 15982
rect 310532 3482 310560 44814
rect 311912 3482 311940 245618
rect 313936 142118 313964 650014
rect 315304 415472 315356 415478
rect 315304 415414 315356 415420
rect 315316 150414 315344 415414
rect 319456 238746 319484 696934
rect 365088 686089 365116 703446
rect 397472 700330 397500 703520
rect 413664 700398 413692 703520
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 399484 700324 399536 700330
rect 399484 700266 399536 700272
rect 365074 686080 365130 686089
rect 365074 686015 365130 686024
rect 364522 685944 364578 685953
rect 364522 685879 364578 685888
rect 364536 678994 364564 685879
rect 364352 678966 364564 678994
rect 364352 676190 364380 678966
rect 364340 676184 364392 676190
rect 364340 676126 364392 676132
rect 364432 666596 364484 666602
rect 364432 666538 364484 666544
rect 364444 659682 364472 666538
rect 364444 659654 364564 659682
rect 364536 654158 364564 659654
rect 364340 654152 364392 654158
rect 364340 654094 364392 654100
rect 364524 654152 364576 654158
rect 364524 654094 364576 654100
rect 364352 644450 364380 654094
rect 364352 644422 364564 644450
rect 364536 634846 364564 644422
rect 364340 634840 364392 634846
rect 364340 634782 364392 634788
rect 364524 634840 364576 634846
rect 364524 634782 364576 634788
rect 364352 625138 364380 634782
rect 364352 625110 364564 625138
rect 364536 615534 364564 625110
rect 364340 615528 364392 615534
rect 364340 615470 364392 615476
rect 364524 615528 364576 615534
rect 364524 615470 364576 615476
rect 364352 605826 364380 615470
rect 364352 605798 364564 605826
rect 364536 596222 364564 605798
rect 364340 596216 364392 596222
rect 364524 596216 364576 596222
rect 364392 596164 364472 596170
rect 364340 596158 364472 596164
rect 364524 596158 364576 596164
rect 364352 596142 364472 596158
rect 364444 596034 364472 596142
rect 364444 596006 364564 596034
rect 364536 591954 364564 596006
rect 364444 591926 364564 591954
rect 364444 589286 364472 591926
rect 364156 589280 364208 589286
rect 364156 589222 364208 589228
rect 364432 589280 364484 589286
rect 364432 589222 364484 589228
rect 364168 579737 364196 589222
rect 364154 579728 364210 579737
rect 329104 579692 329156 579698
rect 364154 579663 364210 579672
rect 364338 579728 364394 579737
rect 364338 579663 364394 579672
rect 329104 579634 329156 579640
rect 322202 267200 322258 267209
rect 322202 267135 322258 267144
rect 319444 238740 319496 238746
rect 319444 238682 319496 238688
rect 316040 160132 316092 160138
rect 316040 160074 316092 160080
rect 315304 150408 315356 150414
rect 315304 150350 315356 150356
rect 313924 142112 313976 142118
rect 313924 142054 313976 142060
rect 313280 103556 313332 103562
rect 313280 103498 313332 103504
rect 306392 3454 307432 3482
rect 307772 3454 308628 3482
rect 309152 3454 309824 3482
rect 310532 3454 311020 3482
rect 311912 3454 312216 3482
rect 307404 480 307432 3454
rect 308600 480 308628 3454
rect 309796 480 309824 3454
rect 310992 480 311020 3454
rect 312188 480 312216 3454
rect 313292 3398 313320 103498
rect 313372 28620 313424 28626
rect 313372 28562 313424 28568
rect 313280 3392 313332 3398
rect 313280 3334 313332 3340
rect 313384 480 313412 28562
rect 315764 9104 315816 9110
rect 315764 9046 315816 9052
rect 314568 3392 314620 3398
rect 314568 3334 314620 3340
rect 314580 480 314608 3334
rect 315776 480 315804 9046
rect 316052 610 316080 160074
rect 318064 87032 318116 87038
rect 318064 86974 318116 86980
rect 318076 47598 318104 86974
rect 318064 47592 318116 47598
rect 318064 47534 318116 47540
rect 318800 24336 318852 24342
rect 318800 24278 318852 24284
rect 318064 9512 318116 9518
rect 318064 9454 318116 9460
rect 316040 604 316092 610
rect 316040 546 316092 552
rect 316960 604 317012 610
rect 316960 546 317012 552
rect 316972 480 317000 546
rect 318076 480 318104 9454
rect 318812 610 318840 24278
rect 320180 21548 320232 21554
rect 320180 21490 320232 21496
rect 320192 626 320220 21490
rect 321560 14680 321612 14686
rect 321560 14622 321612 14628
rect 321572 3398 321600 14622
rect 321652 9376 321704 9382
rect 321652 9318 321704 9324
rect 321560 3392 321612 3398
rect 321560 3334 321612 3340
rect 318800 604 318852 610
rect 318800 546 318852 552
rect 319260 604 319312 610
rect 320192 598 320496 626
rect 319260 546 319312 552
rect 319272 480 319300 546
rect 320468 480 320496 598
rect 321664 480 321692 9318
rect 322216 9110 322244 267135
rect 327080 265328 327132 265334
rect 327080 265270 327132 265276
rect 322296 153264 322348 153270
rect 322296 153206 322348 153212
rect 322308 124166 322336 153206
rect 322296 124160 322348 124166
rect 322296 124102 322348 124108
rect 322940 40860 322992 40866
rect 322940 40802 322992 40808
rect 322204 9104 322256 9110
rect 322204 9046 322256 9052
rect 322848 3392 322900 3398
rect 322848 3334 322900 3340
rect 322860 480 322888 3334
rect 322952 610 322980 40802
rect 324320 22840 324372 22846
rect 324320 22782 324372 22788
rect 324332 610 324360 22782
rect 326436 9036 326488 9042
rect 326436 8978 326488 8984
rect 322940 604 322992 610
rect 322940 546 322992 552
rect 324044 604 324096 610
rect 324044 546 324096 552
rect 324320 604 324372 610
rect 324320 546 324372 552
rect 325240 604 325292 610
rect 325240 546 325292 552
rect 324056 480 324084 546
rect 325252 480 325280 546
rect 326448 480 326476 8978
rect 327092 3482 327120 265270
rect 329116 39982 329144 579634
rect 364352 572642 364380 579663
rect 364352 572614 364472 572642
rect 364444 563122 364472 572614
rect 364444 563094 364564 563122
rect 364536 553450 364564 563094
rect 364524 553444 364576 553450
rect 364524 553386 364576 553392
rect 364524 550656 364576 550662
rect 364524 550598 364576 550604
rect 364536 543862 364564 550598
rect 364524 543856 364576 543862
rect 364524 543798 364576 543804
rect 364616 543788 364668 543794
rect 364616 543730 364668 543736
rect 364628 540977 364656 543730
rect 364430 540968 364486 540977
rect 364430 540903 364486 540912
rect 364614 540968 364670 540977
rect 364614 540903 364670 540912
rect 364444 531350 364472 540903
rect 364432 531344 364484 531350
rect 364432 531286 364484 531292
rect 364708 531344 364760 531350
rect 364708 531286 364760 531292
rect 364720 524550 364748 531286
rect 364708 524544 364760 524550
rect 364708 524486 364760 524492
rect 364616 524408 364668 524414
rect 364616 524350 364668 524356
rect 364628 521665 364656 524350
rect 364430 521656 364486 521665
rect 364430 521591 364486 521600
rect 364614 521656 364670 521665
rect 364614 521591 364670 521600
rect 364444 512038 364472 521591
rect 364432 512032 364484 512038
rect 364432 511974 364484 511980
rect 364708 512032 364760 512038
rect 364708 511974 364760 511980
rect 364720 502382 364748 511974
rect 364524 502376 364576 502382
rect 364246 502344 364302 502353
rect 364246 502279 364302 502288
rect 364522 502344 364524 502353
rect 364708 502376 364760 502382
rect 364576 502344 364578 502353
rect 364708 502318 364760 502324
rect 364522 502279 364578 502288
rect 364260 492697 364288 502279
rect 364246 492688 364302 492697
rect 364246 492623 364302 492632
rect 364430 492688 364486 492697
rect 364430 492623 364486 492632
rect 364444 489954 364472 492623
rect 364444 489926 364564 489954
rect 364536 480282 364564 489926
rect 364340 480276 364392 480282
rect 364340 480218 364392 480224
rect 364524 480276 364576 480282
rect 364524 480218 364576 480224
rect 364352 480162 364380 480218
rect 364352 480134 364472 480162
rect 364444 470642 364472 480134
rect 364444 470614 364564 470642
rect 364536 460970 364564 470614
rect 364340 460964 364392 460970
rect 364340 460906 364392 460912
rect 364524 460964 364576 460970
rect 364524 460906 364576 460912
rect 364352 460850 364380 460906
rect 364352 460822 364472 460850
rect 364444 451330 364472 460822
rect 364444 451302 364564 451330
rect 364536 441658 364564 451302
rect 364340 441652 364392 441658
rect 364340 441594 364392 441600
rect 364524 441652 364576 441658
rect 364524 441594 364576 441600
rect 364352 441538 364380 441594
rect 364352 441510 364472 441538
rect 364444 432018 364472 441510
rect 364444 431990 364564 432018
rect 364536 422346 364564 431990
rect 364340 422340 364392 422346
rect 364340 422282 364392 422288
rect 364524 422340 364576 422346
rect 364524 422282 364576 422288
rect 364352 422226 364380 422282
rect 364352 422198 364472 422226
rect 364444 412706 364472 422198
rect 364444 412678 364564 412706
rect 364536 403034 364564 412678
rect 364340 403028 364392 403034
rect 364340 402970 364392 402976
rect 364524 403028 364576 403034
rect 364524 402970 364576 402976
rect 364352 402914 364380 402970
rect 364352 402886 364472 402914
rect 364444 393394 364472 402886
rect 364444 393366 364564 393394
rect 364536 383722 364564 393366
rect 364340 383716 364392 383722
rect 364340 383658 364392 383664
rect 364524 383716 364576 383722
rect 364524 383658 364576 383664
rect 364352 383602 364380 383658
rect 364352 383574 364472 383602
rect 364444 374082 364472 383574
rect 364444 374054 364564 374082
rect 364536 360262 364564 374054
rect 364524 360256 364576 360262
rect 364524 360198 364576 360204
rect 364524 357536 364576 357542
rect 364524 357478 364576 357484
rect 364536 350554 364564 357478
rect 364352 350526 364564 350554
rect 364352 347750 364380 350526
rect 364340 347744 364392 347750
rect 364340 347686 364392 347692
rect 364432 338156 364484 338162
rect 364432 338098 364484 338104
rect 364444 331242 364472 338098
rect 364444 331214 364564 331242
rect 364536 325718 364564 331214
rect 364340 325712 364392 325718
rect 364340 325654 364392 325660
rect 364524 325712 364576 325718
rect 364524 325654 364576 325660
rect 364352 316010 364380 325654
rect 364352 315982 364564 316010
rect 364536 306406 364564 315982
rect 364340 306400 364392 306406
rect 364340 306342 364392 306348
rect 364524 306400 364576 306406
rect 364524 306342 364576 306348
rect 364352 296698 364380 306342
rect 364352 296670 364564 296698
rect 364536 287094 364564 296670
rect 364340 287088 364392 287094
rect 364340 287030 364392 287036
rect 364524 287088 364576 287094
rect 364524 287030 364576 287036
rect 364352 277386 364380 287030
rect 364352 277358 364564 277386
rect 364536 268433 364564 277358
rect 364522 268424 364578 268433
rect 364522 268359 364578 268368
rect 356702 266520 356758 266529
rect 356702 266455 356758 266464
rect 351920 265668 351972 265674
rect 351920 265610 351972 265616
rect 345020 265600 345072 265606
rect 345020 265542 345072 265548
rect 332600 251252 332652 251258
rect 332600 251194 332652 251200
rect 331220 212560 331272 212566
rect 331220 212502 331272 212508
rect 329104 39976 329156 39982
rect 329104 39918 329156 39924
rect 328460 10328 328512 10334
rect 328460 10270 328512 10276
rect 328472 3482 328500 10270
rect 327092 3454 327672 3482
rect 328472 3454 328868 3482
rect 327644 480 327672 3454
rect 328840 480 328868 3454
rect 330022 3224 330078 3233
rect 330022 3159 330078 3168
rect 330036 480 330064 3159
rect 331232 480 331260 212502
rect 331312 86284 331364 86290
rect 331312 86226 331364 86232
rect 331324 3482 331352 86226
rect 332612 3482 332640 251194
rect 337384 201544 337436 201550
rect 337384 201486 337436 201492
rect 334624 71800 334676 71806
rect 334624 71742 334676 71748
rect 334636 43518 334664 71742
rect 337396 51746 337424 201486
rect 337384 51740 337436 51746
rect 337384 51682 337436 51688
rect 333980 43512 334032 43518
rect 333980 43454 334032 43460
rect 334624 43512 334676 43518
rect 334624 43454 334676 43460
rect 333992 3482 334020 43454
rect 338120 41336 338172 41342
rect 338120 41278 338172 41284
rect 336740 22908 336792 22914
rect 336740 22850 336792 22856
rect 335360 10736 335412 10742
rect 335360 10678 335412 10684
rect 335372 3482 335400 10678
rect 336752 3482 336780 22850
rect 338132 3482 338160 41278
rect 339500 38004 339552 38010
rect 339500 37946 339552 37952
rect 331324 3454 332456 3482
rect 332612 3454 333652 3482
rect 333992 3454 334756 3482
rect 335372 3454 335952 3482
rect 336752 3454 337148 3482
rect 338132 3454 338344 3482
rect 332428 480 332456 3454
rect 333624 480 333652 3454
rect 334728 480 334756 3454
rect 335924 480 335952 3454
rect 337120 480 337148 3454
rect 338316 480 338344 3454
rect 339512 480 339540 37946
rect 340880 35284 340932 35290
rect 340880 35226 340932 35232
rect 340694 4040 340750 4049
rect 340694 3975 340750 3984
rect 340708 480 340736 3975
rect 340892 3482 340920 35226
rect 343640 13184 343692 13190
rect 343640 13126 343692 13132
rect 342260 10668 342312 10674
rect 342260 10610 342312 10616
rect 342272 3482 342300 10610
rect 343652 3482 343680 13126
rect 345032 3482 345060 265542
rect 347780 265124 347832 265130
rect 347780 265066 347832 265072
rect 346400 35216 346452 35222
rect 346400 35158 346452 35164
rect 346412 3482 346440 35158
rect 340892 3454 341932 3482
rect 342272 3454 343128 3482
rect 343652 3454 344324 3482
rect 345032 3454 345520 3482
rect 346412 3454 346716 3482
rect 341904 480 341932 3454
rect 343100 480 343128 3454
rect 344296 480 344324 3454
rect 345492 480 345520 3454
rect 346688 480 346716 3454
rect 347792 3398 347820 265066
rect 347872 117360 347924 117366
rect 347872 117302 347924 117308
rect 347780 3392 347832 3398
rect 347780 3334 347832 3340
rect 347884 480 347912 117302
rect 350540 28416 350592 28422
rect 350540 28358 350592 28364
rect 349160 10464 349212 10470
rect 349160 10406 349212 10412
rect 349172 3482 349200 10406
rect 350552 3482 350580 28358
rect 351932 3482 351960 265610
rect 354680 135312 354732 135318
rect 354680 135254 354732 135260
rect 353300 10532 353352 10538
rect 353300 10474 353352 10480
rect 353312 3482 353340 10474
rect 354692 3482 354720 135254
rect 356060 41064 356112 41070
rect 356060 41006 356112 41012
rect 356072 3482 356100 41006
rect 356152 10396 356204 10402
rect 356152 10338 356204 10344
rect 356164 3942 356192 10338
rect 356716 10334 356744 266455
rect 374000 265736 374052 265742
rect 374000 265678 374052 265684
rect 369860 264036 369912 264042
rect 369860 263978 369912 263984
rect 361580 263968 361632 263974
rect 361580 263910 361632 263916
rect 357440 262948 357492 262954
rect 357440 262890 357492 262896
rect 356704 10328 356756 10334
rect 356704 10270 356756 10276
rect 356152 3936 356204 3942
rect 356152 3878 356204 3884
rect 357348 3936 357400 3942
rect 357348 3878 357400 3884
rect 349172 3454 350304 3482
rect 350552 3454 351408 3482
rect 351932 3454 352604 3482
rect 353312 3454 353800 3482
rect 354692 3454 354996 3482
rect 356072 3454 356192 3482
rect 349068 3392 349120 3398
rect 349068 3334 349120 3340
rect 349080 480 349108 3334
rect 350276 480 350304 3454
rect 351380 480 351408 3454
rect 352576 480 352604 3454
rect 353772 480 353800 3454
rect 354968 480 354996 3454
rect 356164 480 356192 3454
rect 357360 480 357388 3878
rect 357452 3482 357480 262890
rect 358820 74588 358872 74594
rect 358820 74530 358872 74536
rect 358832 3482 358860 74530
rect 360936 9104 360988 9110
rect 360936 9046 360988 9052
rect 357452 3454 358584 3482
rect 358832 3454 359780 3482
rect 358556 480 358584 3454
rect 359752 480 359780 3454
rect 360948 480 360976 9046
rect 361592 3482 361620 263910
rect 368480 263696 368532 263702
rect 368480 263638 368532 263644
rect 367100 258732 367152 258738
rect 367100 258674 367152 258680
rect 364984 187740 365036 187746
rect 364984 187682 365036 187688
rect 362960 43444 363012 43450
rect 362960 43386 363012 43392
rect 362972 3482 363000 43386
rect 364340 10600 364392 10606
rect 364340 10542 364392 10548
rect 364352 3482 364380 10542
rect 364996 10402 365024 187682
rect 365720 41268 365772 41274
rect 365720 41210 365772 41216
rect 364984 10396 365036 10402
rect 364984 10338 365036 10344
rect 361592 3454 362172 3482
rect 362972 3454 363368 3482
rect 364352 3454 364564 3482
rect 362144 480 362172 3454
rect 363340 480 363368 3454
rect 364536 480 364564 3454
rect 365732 3398 365760 41210
rect 365812 6588 365864 6594
rect 365812 6530 365864 6536
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 3210 365852 6530
rect 367112 3482 367140 258674
rect 368492 3482 368520 263638
rect 369872 3482 369900 263978
rect 371884 162920 371936 162926
rect 371884 162862 371936 162868
rect 371240 14544 371292 14550
rect 371240 14486 371292 14492
rect 371252 3482 371280 14486
rect 371896 10470 371924 162862
rect 372620 142180 372672 142186
rect 372620 142122 372672 142128
rect 371884 10464 371936 10470
rect 371884 10406 371936 10412
rect 372632 3482 372660 142122
rect 367112 3454 368060 3482
rect 368492 3454 369256 3482
rect 369872 3454 370452 3482
rect 371252 3454 371648 3482
rect 372632 3454 372844 3482
rect 366916 3392 366968 3398
rect 366916 3334 366968 3340
rect 365732 3182 365852 3210
rect 365732 480 365760 3182
rect 366928 480 366956 3334
rect 368032 480 368060 3454
rect 369228 480 369256 3454
rect 370424 480 370452 3454
rect 371620 480 371648 3454
rect 372816 480 372844 3454
rect 374012 3398 374040 265678
rect 375380 263900 375432 263906
rect 375380 263842 375432 263848
rect 374092 106344 374144 106350
rect 374092 106286 374144 106292
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 1442 374132 106286
rect 375392 3482 375420 263842
rect 390560 263764 390612 263770
rect 390560 263706 390612 263712
rect 385684 216708 385736 216714
rect 385684 216650 385736 216656
rect 380900 41200 380952 41206
rect 380900 41142 380952 41148
rect 376760 40724 376812 40730
rect 376760 40666 376812 40672
rect 376772 3482 376800 40666
rect 379520 36576 379572 36582
rect 379520 36518 379572 36524
rect 378138 29744 378194 29753
rect 378138 29679 378194 29688
rect 378152 3482 378180 29679
rect 379532 3482 379560 36518
rect 380912 3482 380940 41142
rect 383660 40996 383712 41002
rect 383660 40938 383712 40944
rect 382280 10396 382332 10402
rect 382280 10338 382332 10344
rect 382292 3482 382320 10338
rect 383568 6316 383620 6322
rect 383568 6258 383620 6264
rect 375392 3454 376432 3482
rect 376772 3454 377628 3482
rect 378152 3454 378824 3482
rect 379532 3454 380020 3482
rect 380912 3454 381216 3482
rect 382292 3454 382412 3482
rect 375196 3392 375248 3398
rect 375196 3334 375248 3340
rect 374012 1414 374132 1442
rect 374012 480 374040 1414
rect 375208 480 375236 3334
rect 376404 480 376432 3454
rect 377600 480 377628 3454
rect 378796 480 378824 3454
rect 379992 480 380020 3454
rect 381188 480 381216 3454
rect 382384 480 382412 3454
rect 383580 480 383608 6258
rect 383672 3482 383700 40938
rect 385696 11014 385724 216650
rect 389824 95260 389876 95266
rect 389824 95202 389876 95208
rect 386420 45620 386472 45626
rect 386420 45562 386472 45568
rect 385684 11008 385736 11014
rect 385684 10950 385736 10956
rect 385040 10464 385092 10470
rect 385040 10406 385092 10412
rect 385052 3482 385080 10406
rect 386432 3482 386460 45562
rect 389180 11008 389232 11014
rect 389180 10950 389232 10956
rect 388260 6724 388312 6730
rect 388260 6666 388312 6672
rect 383672 3454 384712 3482
rect 385052 3454 385908 3482
rect 386432 3454 387104 3482
rect 384684 480 384712 3454
rect 385880 480 385908 3454
rect 387076 480 387104 3454
rect 388272 480 388300 6666
rect 389192 3482 389220 10950
rect 389836 10402 389864 95202
rect 389824 10396 389876 10402
rect 389824 10338 389876 10344
rect 390572 3482 390600 263706
rect 396080 238060 396132 238066
rect 396080 238002 396132 238008
rect 390652 39364 390704 39370
rect 390652 39306 390704 39312
rect 390664 3942 390692 39306
rect 391940 25560 391992 25566
rect 391940 25502 391992 25508
rect 390652 3936 390704 3942
rect 390652 3878 390704 3884
rect 391848 3936 391900 3942
rect 391848 3878 391900 3884
rect 389192 3454 389496 3482
rect 390572 3454 390692 3482
rect 389468 480 389496 3454
rect 390664 480 390692 3454
rect 391860 480 391888 3878
rect 391952 3482 391980 25502
rect 393318 21312 393374 21321
rect 393318 21247 393374 21256
rect 391952 3454 393084 3482
rect 393056 480 393084 3454
rect 393332 610 393360 21247
rect 395436 7880 395488 7886
rect 395436 7822 395488 7828
rect 393320 604 393372 610
rect 393320 546 393372 552
rect 394240 604 394292 610
rect 394240 546 394292 552
rect 394252 480 394280 546
rect 395448 480 395476 7822
rect 396092 610 396120 238002
rect 399496 42537 399524 700266
rect 429856 688634 429884 703520
rect 429384 688628 429436 688634
rect 429384 688570 429436 688576
rect 429844 688628 429896 688634
rect 429844 688570 429896 688576
rect 429396 685930 429424 688570
rect 429304 685902 429424 685930
rect 429304 684486 429332 685902
rect 429292 684480 429344 684486
rect 429292 684422 429344 684428
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 429672 659682 429700 666538
rect 429488 659654 429700 659682
rect 429488 647290 429516 659654
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 429396 640422 429424 647226
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 429488 630698 429516 640358
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 429304 630578 429332 630634
rect 429304 630550 429424 630578
rect 429396 621058 429424 630550
rect 429396 621030 429516 621058
rect 429488 611386 429516 621030
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 429304 611266 429332 611322
rect 429304 611238 429424 611266
rect 429396 608598 429424 611238
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 429580 598942 429608 601666
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 429660 589348 429712 589354
rect 429660 589290 429712 589296
rect 429672 582486 429700 589290
rect 429660 582480 429712 582486
rect 429660 582422 429712 582428
rect 429568 582344 429620 582350
rect 429568 582286 429620 582292
rect 429580 572642 429608 582286
rect 429396 572614 429608 572642
rect 429396 569922 429424 572614
rect 429304 569894 429424 569922
rect 429304 563174 429332 569894
rect 429292 563168 429344 563174
rect 429292 563110 429344 563116
rect 429292 563032 429344 563038
rect 429292 562974 429344 562980
rect 429304 560250 429332 562974
rect 429292 560244 429344 560250
rect 429292 560186 429344 560192
rect 424874 556472 424930 556481
rect 424874 556407 424930 556416
rect 425058 556472 425114 556481
rect 425058 556407 425114 556416
rect 424888 556374 424916 556407
rect 415400 556368 415452 556374
rect 415398 556336 415400 556345
rect 424876 556368 424928 556374
rect 415452 556336 415454 556345
rect 424876 556310 424928 556316
rect 415398 556271 415454 556280
rect 425072 555937 425100 556407
rect 425058 555928 425114 555937
rect 425058 555863 425114 555872
rect 429476 550656 429528 550662
rect 429476 550598 429528 550604
rect 429488 543658 429516 550598
rect 429292 543652 429344 543658
rect 429292 543594 429344 543600
rect 429476 543652 429528 543658
rect 429476 543594 429528 543600
rect 429304 534070 429332 543594
rect 429292 534064 429344 534070
rect 429292 534006 429344 534012
rect 429476 534064 429528 534070
rect 429476 534006 429528 534012
rect 429488 524482 429516 534006
rect 429476 524476 429528 524482
rect 429476 524418 429528 524424
rect 429568 524408 429620 524414
rect 429568 524350 429620 524356
rect 429580 521665 429608 524350
rect 429382 521656 429438 521665
rect 429382 521591 429438 521600
rect 429566 521656 429622 521665
rect 429566 521591 429622 521600
rect 429396 512038 429424 521591
rect 429384 512032 429436 512038
rect 429384 511974 429436 511980
rect 429660 512032 429712 512038
rect 429660 511974 429712 511980
rect 429672 502382 429700 511974
rect 429476 502376 429528 502382
rect 429198 502344 429254 502353
rect 429198 502279 429254 502288
rect 429474 502344 429476 502353
rect 429660 502376 429712 502382
rect 429528 502344 429530 502353
rect 429660 502318 429712 502324
rect 429474 502279 429530 502288
rect 429212 492697 429240 502279
rect 429198 492688 429254 492697
rect 429198 492623 429254 492632
rect 429382 492688 429438 492697
rect 429382 492623 429384 492632
rect 429436 492623 429438 492632
rect 429384 492594 429436 492600
rect 429384 485784 429436 485790
rect 429384 485726 429436 485732
rect 429396 483018 429424 485726
rect 429396 482990 429516 483018
rect 429488 476134 429516 482990
rect 429292 476128 429344 476134
rect 429476 476128 429528 476134
rect 429344 476076 429424 476082
rect 429292 476070 429424 476076
rect 429476 476070 429528 476076
rect 429304 476054 429424 476070
rect 429396 473346 429424 476054
rect 429384 473340 429436 473346
rect 429384 473282 429436 473288
rect 429384 466404 429436 466410
rect 429384 466346 429436 466352
rect 429396 463706 429424 466346
rect 429396 463678 429516 463706
rect 429488 454073 429516 463678
rect 429198 454064 429254 454073
rect 429198 453999 429254 454008
rect 429474 454064 429530 454073
rect 429474 453999 429530 454008
rect 429212 447166 429240 453999
rect 429200 447160 429252 447166
rect 429200 447102 429252 447108
rect 429292 447092 429344 447098
rect 429292 447034 429344 447040
rect 429304 444378 429332 447034
rect 429016 444372 429068 444378
rect 429016 444314 429068 444320
rect 429292 444372 429344 444378
rect 429292 444314 429344 444320
rect 429028 434761 429056 444314
rect 429014 434752 429070 434761
rect 429014 434687 429070 434696
rect 429198 434752 429254 434761
rect 429198 434687 429254 434696
rect 429212 427854 429240 434687
rect 429200 427848 429252 427854
rect 429200 427790 429252 427796
rect 429292 427780 429344 427786
rect 429292 427722 429344 427728
rect 429304 425066 429332 427722
rect 429016 425060 429068 425066
rect 429016 425002 429068 425008
rect 429292 425060 429344 425066
rect 429292 425002 429344 425008
rect 429028 415449 429056 425002
rect 429014 415440 429070 415449
rect 429014 415375 429070 415384
rect 429198 415440 429254 415449
rect 429198 415375 429254 415384
rect 429212 408542 429240 415375
rect 429200 408536 429252 408542
rect 429200 408478 429252 408484
rect 429292 408400 429344 408406
rect 429292 408342 429344 408348
rect 429304 405686 429332 408342
rect 429292 405680 429344 405686
rect 429292 405622 429344 405628
rect 429292 398812 429344 398818
rect 429292 398754 429344 398760
rect 429304 389230 429332 398754
rect 429292 389224 429344 389230
rect 429292 389166 429344 389172
rect 429292 389088 429344 389094
rect 429292 389030 429344 389036
rect 429304 379506 429332 389030
rect 429292 379500 429344 379506
rect 429292 379442 429344 379448
rect 429476 379500 429528 379506
rect 429476 379442 429528 379448
rect 429488 371906 429516 379442
rect 429488 371878 429608 371906
rect 429580 357542 429608 371878
rect 429568 357536 429620 357542
rect 429568 357478 429620 357484
rect 429568 353388 429620 353394
rect 429568 353330 429620 353336
rect 429580 353274 429608 353330
rect 429580 353258 429700 353274
rect 429580 353252 429712 353258
rect 429580 353246 429660 353252
rect 429660 353194 429712 353200
rect 429660 340808 429712 340814
rect 429660 340750 429712 340756
rect 429672 331514 429700 340750
rect 429580 331486 429700 331514
rect 429580 325718 429608 331486
rect 429476 325712 429528 325718
rect 429476 325654 429528 325660
rect 429568 325712 429620 325718
rect 429568 325654 429620 325660
rect 429488 318850 429516 325654
rect 429384 318844 429436 318850
rect 429384 318786 429436 318792
rect 429476 318844 429528 318850
rect 429476 318786 429528 318792
rect 429396 311982 429424 318786
rect 429384 311976 429436 311982
rect 429384 311918 429436 311924
rect 429476 311976 429528 311982
rect 429476 311918 429528 311924
rect 429488 302258 429516 311918
rect 429292 302252 429344 302258
rect 429292 302194 429344 302200
rect 429476 302252 429528 302258
rect 429476 302194 429528 302200
rect 429304 302138 429332 302194
rect 429304 302110 429424 302138
rect 429396 292482 429424 302110
rect 429396 292454 429516 292482
rect 429488 289814 429516 292454
rect 429476 289808 429528 289814
rect 429476 289750 429528 289756
rect 429568 280220 429620 280226
rect 429568 280162 429620 280168
rect 429580 274922 429608 280162
rect 429384 274916 429436 274922
rect 429384 274858 429436 274864
rect 429568 274916 429620 274922
rect 429568 274858 429620 274864
rect 429396 270502 429424 274858
rect 462332 272542 462360 703520
rect 478524 700330 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700324 478564 700330
rect 478512 700266 478564 700272
rect 494900 686089 494928 703446
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 494242 685944 494298 685953
rect 494242 685879 494298 685888
rect 494256 678994 494284 685879
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 494164 659682 494192 666538
rect 494164 659654 494284 659682
rect 494256 654158 494284 659654
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 494072 644450 494100 654094
rect 494072 644422 494284 644450
rect 494256 634846 494284 644422
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 494072 625138 494100 634782
rect 494072 625110 494284 625138
rect 494256 615534 494284 625110
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 494072 605826 494100 615470
rect 494072 605798 494284 605826
rect 494256 596222 494284 605798
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 494256 591954 494284 596006
rect 494164 591926 494284 591954
rect 494164 589286 494192 591926
rect 493876 589280 493928 589286
rect 493876 589222 493928 589228
rect 494152 589280 494204 589286
rect 494152 589222 494204 589228
rect 493888 579737 493916 589222
rect 493874 579728 493930 579737
rect 493874 579663 493930 579672
rect 494058 579728 494114 579737
rect 494058 579663 494114 579672
rect 494072 572642 494100 579663
rect 494072 572614 494192 572642
rect 494164 563122 494192 572614
rect 494164 563094 494284 563122
rect 494256 553450 494284 563094
rect 521658 556472 521714 556481
rect 521658 556407 521660 556416
rect 521712 556407 521714 556416
rect 521660 556378 521712 556384
rect 494244 553444 494296 553450
rect 494244 553386 494296 553392
rect 494244 550656 494296 550662
rect 494244 550598 494296 550604
rect 494256 543862 494284 550598
rect 494244 543856 494296 543862
rect 494244 543798 494296 543804
rect 494336 543788 494388 543794
rect 494336 543730 494388 543736
rect 494348 540977 494376 543730
rect 494150 540968 494206 540977
rect 494150 540903 494206 540912
rect 494334 540968 494390 540977
rect 494334 540903 494390 540912
rect 494164 531350 494192 540903
rect 494152 531344 494204 531350
rect 494152 531286 494204 531292
rect 494428 531344 494480 531350
rect 494428 531286 494480 531292
rect 494440 524550 494468 531286
rect 494428 524544 494480 524550
rect 494428 524486 494480 524492
rect 494336 524408 494388 524414
rect 494336 524350 494388 524356
rect 494348 521665 494376 524350
rect 494150 521656 494206 521665
rect 494150 521591 494206 521600
rect 494334 521656 494390 521665
rect 494334 521591 494390 521600
rect 494164 512038 494192 521591
rect 494152 512032 494204 512038
rect 494152 511974 494204 511980
rect 494428 512032 494480 512038
rect 494428 511974 494480 511980
rect 494440 502382 494468 511974
rect 494244 502376 494296 502382
rect 493966 502344 494022 502353
rect 493966 502279 494022 502288
rect 494242 502344 494244 502353
rect 494428 502376 494480 502382
rect 494296 502344 494298 502353
rect 494428 502318 494480 502324
rect 494242 502279 494298 502288
rect 493980 492697 494008 502279
rect 493966 492688 494022 492697
rect 493966 492623 494022 492632
rect 494150 492688 494206 492697
rect 494150 492623 494206 492632
rect 494164 489954 494192 492623
rect 494164 489926 494284 489954
rect 494256 480282 494284 489926
rect 494060 480276 494112 480282
rect 494060 480218 494112 480224
rect 494244 480276 494296 480282
rect 494244 480218 494296 480224
rect 494072 480162 494100 480218
rect 494072 480134 494192 480162
rect 494164 470642 494192 480134
rect 494164 470614 494284 470642
rect 494256 460970 494284 470614
rect 494060 460964 494112 460970
rect 494060 460906 494112 460912
rect 494244 460964 494296 460970
rect 494244 460906 494296 460912
rect 494072 460850 494100 460906
rect 494072 460822 494192 460850
rect 494164 451330 494192 460822
rect 494164 451302 494284 451330
rect 494256 441658 494284 451302
rect 494060 441652 494112 441658
rect 494060 441594 494112 441600
rect 494244 441652 494296 441658
rect 494244 441594 494296 441600
rect 494072 441538 494100 441594
rect 494072 441510 494192 441538
rect 494164 432018 494192 441510
rect 494164 431990 494284 432018
rect 494256 422346 494284 431990
rect 494060 422340 494112 422346
rect 494060 422282 494112 422288
rect 494244 422340 494296 422346
rect 494244 422282 494296 422288
rect 494072 422226 494100 422282
rect 494072 422198 494192 422226
rect 494164 412706 494192 422198
rect 494164 412678 494284 412706
rect 494256 403034 494284 412678
rect 494060 403028 494112 403034
rect 494060 402970 494112 402976
rect 494244 403028 494296 403034
rect 494244 402970 494296 402976
rect 494072 402914 494100 402970
rect 494072 402886 494192 402914
rect 494164 393394 494192 402886
rect 494164 393366 494284 393394
rect 494256 383722 494284 393366
rect 494060 383716 494112 383722
rect 494060 383658 494112 383664
rect 494244 383716 494296 383722
rect 494244 383658 494296 383664
rect 494072 383602 494100 383658
rect 494072 383574 494192 383602
rect 494164 374082 494192 383574
rect 494164 374054 494284 374082
rect 494256 360262 494284 374054
rect 494244 360256 494296 360262
rect 494244 360198 494296 360204
rect 494244 357536 494296 357542
rect 494244 357478 494296 357484
rect 494256 350554 494284 357478
rect 494072 350526 494284 350554
rect 494072 347750 494100 350526
rect 494060 347744 494112 347750
rect 494060 347686 494112 347692
rect 494152 338156 494204 338162
rect 494152 338098 494204 338104
rect 494164 331242 494192 338098
rect 494164 331214 494284 331242
rect 494256 325718 494284 331214
rect 494060 325712 494112 325718
rect 494060 325654 494112 325660
rect 494244 325712 494296 325718
rect 494244 325654 494296 325660
rect 494072 316010 494100 325654
rect 494072 315982 494284 316010
rect 494256 306406 494284 315982
rect 494060 306400 494112 306406
rect 494060 306342 494112 306348
rect 494244 306400 494296 306406
rect 494244 306342 494296 306348
rect 494072 296698 494100 306342
rect 494072 296670 494284 296698
rect 494256 287094 494284 296670
rect 494060 287088 494112 287094
rect 494060 287030 494112 287036
rect 494244 287088 494296 287094
rect 494244 287030 494296 287036
rect 494072 282198 494100 287030
rect 494060 282192 494112 282198
rect 494060 282134 494112 282140
rect 462320 272536 462372 272542
rect 462320 272478 462372 272484
rect 527192 271182 527220 703520
rect 543476 703474 543504 703520
rect 543476 703446 543596 703474
rect 533344 700324 533396 700330
rect 533344 700266 533396 700272
rect 529296 556436 529348 556442
rect 529296 556378 529348 556384
rect 529308 556209 529336 556378
rect 529294 556200 529350 556209
rect 529294 556135 529350 556144
rect 527180 271176 527232 271182
rect 527180 271118 527232 271124
rect 443000 270700 443052 270706
rect 443000 270642 443052 270648
rect 429384 270496 429436 270502
rect 429384 270438 429436 270444
rect 412640 269544 412692 269550
rect 412640 269486 412692 269492
rect 408500 268320 408552 268326
rect 408500 268262 408552 268268
rect 407762 267880 407818 267889
rect 407762 267815 407818 267824
rect 402980 256012 403032 256018
rect 402980 255954 403032 255960
rect 400220 243568 400272 243574
rect 400220 243510 400272 243516
rect 399482 42528 399538 42537
rect 399482 42463 399538 42472
rect 397826 9072 397882 9081
rect 397826 9007 397882 9016
rect 396080 604 396132 610
rect 396080 546 396132 552
rect 396632 604 396684 610
rect 396632 546 396684 552
rect 396644 480 396672 546
rect 397840 480 397868 9007
rect 399024 7676 399076 7682
rect 399024 7618 399076 7624
rect 399036 480 399064 7618
rect 400232 480 400260 243510
rect 401600 24268 401652 24274
rect 401600 24210 401652 24216
rect 401322 6896 401378 6905
rect 401322 6831 401378 6840
rect 401336 480 401364 6831
rect 401612 610 401640 24210
rect 402992 3346 403020 255954
rect 403624 78736 403676 78742
rect 403624 78678 403676 78684
rect 403636 4078 403664 78678
rect 407776 64870 407804 267815
rect 407764 64864 407816 64870
rect 407764 64806 407816 64812
rect 405740 41132 405792 41138
rect 405740 41074 405792 41080
rect 404912 6656 404964 6662
rect 404912 6598 404964 6604
rect 403624 4072 403676 4078
rect 403624 4014 403676 4020
rect 402992 3318 403756 3346
rect 401600 604 401652 610
rect 401600 546 401652 552
rect 402520 604 402572 610
rect 402520 546 402572 552
rect 402532 480 402560 546
rect 403728 480 403756 3318
rect 404924 480 404952 6598
rect 405752 3346 405780 41074
rect 407764 40792 407816 40798
rect 407764 40734 407816 40740
rect 407120 10396 407172 10402
rect 407120 10338 407172 10344
rect 407132 3346 407160 10338
rect 407776 4010 407804 40734
rect 407764 4004 407816 4010
rect 407764 3946 407816 3952
rect 408512 3942 408540 268262
rect 411260 107704 411312 107710
rect 411260 107646 411312 107652
rect 409144 98048 409196 98054
rect 409144 97990 409196 97996
rect 408592 11892 408644 11898
rect 408592 11834 408644 11840
rect 408500 3936 408552 3942
rect 408500 3878 408552 3884
rect 408604 3482 408632 11834
rect 409156 11014 409184 97990
rect 409144 11008 409196 11014
rect 409144 10950 409196 10956
rect 409880 11008 409932 11014
rect 409880 10950 409932 10956
rect 409696 3936 409748 3942
rect 409696 3878 409748 3884
rect 408512 3454 408632 3482
rect 405752 3318 406148 3346
rect 407132 3318 407344 3346
rect 406120 480 406148 3318
rect 407316 480 407344 3318
rect 408512 480 408540 3454
rect 409708 480 409736 3878
rect 409892 3346 409920 10950
rect 411272 3346 411300 107646
rect 409892 3318 410932 3346
rect 411272 3318 412128 3346
rect 410904 480 410932 3318
rect 412100 480 412128 3318
rect 412652 610 412680 269486
rect 418160 269476 418212 269482
rect 418160 269418 418212 269424
rect 416872 269408 416924 269414
rect 416872 269350 416924 269356
rect 415398 33824 415454 33833
rect 415398 33759 415454 33768
rect 414020 15972 414072 15978
rect 414020 15914 414072 15920
rect 414032 626 414060 15914
rect 412640 604 412692 610
rect 412640 546 412692 552
rect 413284 604 413336 610
rect 414032 598 414520 626
rect 415412 610 415440 33759
rect 413284 546 413336 552
rect 413296 480 413324 546
rect 414492 480 414520 598
rect 415400 604 415452 610
rect 415400 546 415452 552
rect 415676 604 415728 610
rect 415676 546 415728 552
rect 415688 480 415716 546
rect 416884 480 416912 269350
rect 417976 3868 418028 3874
rect 417976 3810 418028 3816
rect 417988 480 418016 3810
rect 418172 610 418200 269418
rect 419540 269272 419592 269278
rect 419540 269214 419592 269220
rect 419552 610 419580 269214
rect 436100 268252 436152 268258
rect 436100 268194 436152 268200
rect 435364 265192 435416 265198
rect 435364 265134 435416 265140
rect 429384 263560 429436 263566
rect 429384 263502 429436 263508
rect 429396 260846 429424 263502
rect 429384 260840 429436 260846
rect 429384 260782 429436 260788
rect 429568 253972 429620 253978
rect 429568 253914 429620 253920
rect 429580 244202 429608 253914
rect 429396 244174 429608 244202
rect 429396 241482 429424 244174
rect 429304 241454 429424 241482
rect 429304 234734 429332 241454
rect 429292 234728 429344 234734
rect 429292 234670 429344 234676
rect 429292 234592 429344 234598
rect 429292 234534 429344 234540
rect 429304 231810 429332 234534
rect 429292 231804 429344 231810
rect 429292 231746 429344 231752
rect 429476 222216 429528 222222
rect 429476 222158 429528 222164
rect 429488 215218 429516 222158
rect 429292 215212 429344 215218
rect 429292 215154 429344 215160
rect 429476 215212 429528 215218
rect 429476 215154 429528 215160
rect 429304 205630 429332 215154
rect 429292 205624 429344 205630
rect 429292 205566 429344 205572
rect 429476 205624 429528 205630
rect 429476 205566 429528 205572
rect 429488 202842 429516 205566
rect 429476 202836 429528 202842
rect 429476 202778 429528 202784
rect 430580 198756 430632 198762
rect 430580 198698 430632 198704
rect 429568 193316 429620 193322
rect 429568 193258 429620 193264
rect 429580 186266 429608 193258
rect 429488 186238 429608 186266
rect 429488 183530 429516 186238
rect 429476 183524 429528 183530
rect 429476 183466 429528 183472
rect 429568 174004 429620 174010
rect 429568 173946 429620 173952
rect 429580 166954 429608 173946
rect 429396 166926 429608 166954
rect 429396 164218 429424 166926
rect 429384 164212 429436 164218
rect 429384 164154 429436 164160
rect 422944 157412 422996 157418
rect 422944 157354 422996 157360
rect 422956 144906 422984 157354
rect 429384 157344 429436 157350
rect 429384 157286 429436 157292
rect 429396 154578 429424 157286
rect 429396 154550 429516 154578
rect 429488 147694 429516 154550
rect 429292 147688 429344 147694
rect 429476 147688 429528 147694
rect 429344 147636 429424 147642
rect 429292 147630 429424 147636
rect 429476 147630 429528 147636
rect 429304 147614 429424 147630
rect 429396 144906 429424 147614
rect 422944 144900 422996 144906
rect 422944 144842 422996 144848
rect 429384 144900 429436 144906
rect 429384 144842 429436 144848
rect 429384 137964 429436 137970
rect 429384 137906 429436 137912
rect 426440 136672 426492 136678
rect 426440 136614 426492 136620
rect 423680 109064 423732 109070
rect 423680 109006 423732 109012
rect 422760 6384 422812 6390
rect 422760 6326 422812 6332
rect 421564 3800 421616 3806
rect 421564 3742 421616 3748
rect 418160 604 418212 610
rect 418160 546 418212 552
rect 419172 604 419224 610
rect 419172 546 419224 552
rect 419540 604 419592 610
rect 419540 546 419592 552
rect 420368 604 420420 610
rect 420368 546 420420 552
rect 419184 480 419212 546
rect 420380 480 420408 546
rect 421576 480 421604 3742
rect 422772 480 422800 6326
rect 423692 3482 423720 109006
rect 425152 37936 425204 37942
rect 425152 37878 425204 37884
rect 425060 3664 425112 3670
rect 425060 3606 425112 3612
rect 423692 3454 423996 3482
rect 423968 480 423996 3454
rect 425072 3346 425100 3606
rect 425164 3534 425192 37878
rect 425152 3528 425204 3534
rect 425152 3470 425204 3476
rect 426348 3528 426400 3534
rect 426348 3470 426400 3476
rect 426452 3482 426480 136614
rect 429396 135266 429424 137906
rect 429396 135238 429516 135266
rect 429488 128382 429516 135238
rect 429292 128376 429344 128382
rect 429292 128318 429344 128324
rect 429476 128376 429528 128382
rect 429476 128318 429528 128324
rect 429304 125594 429332 128318
rect 429292 125588 429344 125594
rect 429292 125530 429344 125536
rect 429292 116000 429344 116006
rect 429292 115942 429344 115948
rect 429304 109018 429332 115942
rect 429304 108990 429516 109018
rect 429488 101402 429516 108990
rect 429396 101374 429516 101402
rect 429396 96626 429424 101374
rect 429108 96620 429160 96626
rect 429108 96562 429160 96568
rect 429384 96620 429436 96626
rect 429384 96562 429436 96568
rect 429120 87009 429148 96562
rect 429106 87000 429162 87009
rect 429106 86935 429162 86944
rect 429290 87000 429346 87009
rect 429290 86935 429346 86944
rect 429304 80102 429332 86935
rect 429292 80096 429344 80102
rect 429292 80038 429344 80044
rect 429384 79960 429436 79966
rect 429384 79902 429436 79908
rect 429396 70530 429424 79902
rect 429396 70502 429516 70530
rect 429488 70258 429516 70502
rect 429304 70230 429516 70258
rect 429304 67561 429332 70230
rect 429290 67552 429346 67561
rect 429290 67487 429346 67496
rect 429566 67552 429622 67561
rect 429566 67487 429622 67496
rect 429580 60654 429608 67487
rect 429384 60648 429436 60654
rect 429384 60590 429436 60596
rect 429568 60648 429620 60654
rect 429568 60590 429620 60596
rect 429396 42838 429424 60590
rect 429384 42832 429436 42838
rect 429384 42774 429436 42780
rect 429198 35184 429254 35193
rect 429198 35119 429254 35128
rect 429212 3482 429240 35119
rect 430592 3482 430620 198698
rect 433340 111852 433392 111858
rect 433340 111794 433392 111800
rect 432328 3936 432380 3942
rect 432328 3878 432380 3884
rect 425072 3318 425192 3346
rect 425164 480 425192 3318
rect 426360 480 426388 3470
rect 426452 3454 427584 3482
rect 429212 3454 429976 3482
rect 430592 3454 431172 3482
rect 427556 480 427584 3454
rect 428740 3392 428792 3398
rect 428740 3334 428792 3340
rect 428752 480 428780 3334
rect 429948 480 429976 3454
rect 431144 480 431172 3454
rect 432340 480 432368 3878
rect 433352 3534 433380 111794
rect 433432 85604 433484 85610
rect 433432 85546 433484 85552
rect 433340 3528 433392 3534
rect 433340 3470 433392 3476
rect 433444 3482 433472 85546
rect 435376 3534 435404 265134
rect 435824 4004 435876 4010
rect 435824 3946 435876 3952
rect 434628 3528 434680 3534
rect 433444 3454 433564 3482
rect 434628 3470 434680 3476
rect 435364 3528 435416 3534
rect 435364 3470 435416 3476
rect 433536 480 433564 3454
rect 434640 480 434668 3470
rect 435836 480 435864 3946
rect 436112 3482 436140 268194
rect 437480 265260 437532 265266
rect 437480 265202 437532 265208
rect 437492 3482 437520 265202
rect 441620 40928 441672 40934
rect 441620 40870 441672 40876
rect 438860 31068 438912 31074
rect 438860 31010 438912 31016
rect 438872 3482 438900 31010
rect 440608 6180 440660 6186
rect 440608 6122 440660 6128
rect 436112 3454 437060 3482
rect 437492 3454 438256 3482
rect 438872 3454 439452 3482
rect 437032 480 437060 3454
rect 438228 480 438256 3454
rect 439424 480 439452 3454
rect 440620 480 440648 6122
rect 441632 3482 441660 40870
rect 441632 3454 441844 3482
rect 441816 480 441844 3454
rect 443012 3398 443040 270642
rect 458180 270632 458232 270638
rect 458180 270574 458232 270580
rect 451280 263832 451332 263838
rect 451280 263774 451332 263780
rect 445760 262880 445812 262886
rect 445760 262822 445812 262828
rect 443092 17400 443144 17406
rect 443092 17342 443144 17348
rect 443000 3392 443052 3398
rect 443000 3334 443052 3340
rect 443104 1442 443132 17342
rect 444380 11756 444432 11762
rect 444380 11698 444432 11704
rect 444392 3482 444420 11698
rect 445772 3482 445800 262822
rect 447140 171148 447192 171154
rect 447140 171090 447192 171096
rect 447152 3482 447180 171090
rect 448520 33856 448572 33862
rect 448520 33798 448572 33804
rect 448532 3482 448560 33798
rect 450174 3768 450230 3777
rect 450174 3703 450230 3712
rect 444392 3454 445432 3482
rect 445772 3454 446628 3482
rect 447152 3454 447824 3482
rect 448532 3454 449020 3482
rect 444196 3392 444248 3398
rect 444196 3334 444248 3340
rect 443012 1414 443132 1442
rect 443012 480 443040 1414
rect 444208 480 444236 3334
rect 445404 480 445432 3454
rect 446600 480 446628 3454
rect 447796 480 447824 3454
rect 448992 480 449020 3454
rect 450188 480 450216 3703
rect 451292 480 451320 263774
rect 451372 261588 451424 261594
rect 451372 261530 451424 261536
rect 451384 3482 451412 261530
rect 455420 260228 455472 260234
rect 455420 260170 455472 260176
rect 454866 8936 454922 8945
rect 454866 8871 454922 8880
rect 453672 4888 453724 4894
rect 453672 4830 453724 4836
rect 451384 3454 452516 3482
rect 452488 480 452516 3454
rect 453684 480 453712 4830
rect 454880 480 454908 8871
rect 455432 3482 455460 260170
rect 457258 3632 457314 3641
rect 457258 3567 457314 3576
rect 455432 3454 456104 3482
rect 456076 480 456104 3454
rect 457272 480 457300 3567
rect 458192 3482 458220 270574
rect 476120 270564 476172 270570
rect 476120 270506 476172 270512
rect 460940 270020 460992 270026
rect 460940 269962 460992 269968
rect 459560 261520 459612 261526
rect 459560 261462 459612 261468
rect 459572 3482 459600 261462
rect 459652 50380 459704 50386
rect 459652 50322 459704 50328
rect 459664 3670 459692 50322
rect 459652 3664 459704 3670
rect 459652 3606 459704 3612
rect 460848 3664 460900 3670
rect 460848 3606 460900 3612
rect 458192 3454 458496 3482
rect 459572 3454 459692 3482
rect 458468 480 458496 3454
rect 459664 480 459692 3454
rect 460860 480 460888 3606
rect 460952 3482 460980 269962
rect 465080 269340 465132 269346
rect 465080 269282 465132 269288
rect 462320 211200 462372 211206
rect 462320 211142 462372 211148
rect 462332 3482 462360 211142
rect 463700 10328 463752 10334
rect 463700 10270 463752 10276
rect 463712 3482 463740 10270
rect 465092 3482 465120 269282
rect 467840 257372 467892 257378
rect 467840 257314 467892 257320
rect 467104 226364 467156 226370
rect 467104 226306 467156 226312
rect 466460 22772 466512 22778
rect 466460 22714 466512 22720
rect 466472 3482 466500 22714
rect 467116 3670 467144 226306
rect 467104 3664 467156 3670
rect 467104 3606 467156 3612
rect 460952 3454 462084 3482
rect 462332 3454 463280 3482
rect 463712 3454 464476 3482
rect 465092 3454 465672 3482
rect 466472 3454 466868 3482
rect 462056 480 462084 3454
rect 463252 480 463280 3454
rect 464448 480 464476 3454
rect 465644 480 465672 3454
rect 466840 480 466868 3454
rect 467852 1578 467880 257314
rect 469220 89752 469272 89758
rect 469220 89694 469272 89700
rect 467932 24132 467984 24138
rect 467932 24074 467984 24080
rect 467944 3398 467972 24074
rect 469232 3482 469260 89694
rect 473358 25664 473414 25673
rect 473358 25599 473414 25608
rect 471978 25528 472034 25537
rect 471978 25463 472034 25472
rect 471520 3596 471572 3602
rect 471520 3538 471572 3544
rect 469232 3454 470364 3482
rect 467932 3392 467984 3398
rect 467932 3334 467984 3340
rect 469128 3392 469180 3398
rect 469128 3334 469180 3340
rect 467852 1550 467972 1578
rect 467944 480 467972 1550
rect 469140 480 469168 3334
rect 470336 480 470364 3454
rect 471532 480 471560 3538
rect 471992 3482 472020 25463
rect 473372 3482 473400 25599
rect 475108 3732 475160 3738
rect 475108 3674 475160 3680
rect 471992 3454 472756 3482
rect 473372 3454 473952 3482
rect 472728 480 472756 3454
rect 473924 480 473952 3454
rect 475120 480 475148 3674
rect 476132 3482 476160 270506
rect 520280 269952 520332 269958
rect 520280 269894 520332 269900
rect 487158 269240 487214 269249
rect 487158 269175 487214 269184
rect 482284 265872 482336 265878
rect 482284 265814 482336 265820
rect 478880 207052 478932 207058
rect 478880 206994 478932 207000
rect 477500 173936 477552 173942
rect 477500 173878 477552 173884
rect 476132 3454 476344 3482
rect 476316 480 476344 3454
rect 477512 480 477540 173878
rect 478696 9240 478748 9246
rect 478696 9182 478748 9188
rect 478708 480 478736 9182
rect 478892 3482 478920 206994
rect 480258 29608 480314 29617
rect 480258 29543 480314 29552
rect 480272 3482 480300 29543
rect 482296 5114 482324 265814
rect 485780 260160 485832 260166
rect 485780 260102 485832 260108
rect 483020 32428 483072 32434
rect 483020 32370 483072 32376
rect 482296 5086 482416 5114
rect 478892 3454 479932 3482
rect 480272 3454 481128 3482
rect 482388 3466 482416 5086
rect 483032 3482 483060 32370
rect 484400 28348 484452 28354
rect 484400 28290 484452 28296
rect 484412 3482 484440 28290
rect 479904 480 479932 3454
rect 481100 480 481128 3454
rect 482284 3460 482336 3466
rect 482284 3402 482336 3408
rect 482376 3460 482428 3466
rect 483032 3454 483520 3482
rect 484412 3454 484624 3482
rect 482376 3402 482428 3408
rect 482296 480 482324 3402
rect 483492 480 483520 3454
rect 484596 480 484624 3454
rect 485792 480 485820 260102
rect 486974 3496 487030 3505
rect 487172 3482 487200 269175
rect 518900 268048 518952 268054
rect 518900 267990 518952 267996
rect 494058 266656 494114 266665
rect 494058 266591 494114 266600
rect 492680 264240 492732 264246
rect 492680 264182 492732 264188
rect 491300 120148 491352 120154
rect 491300 120090 491352 120096
rect 488540 18624 488592 18630
rect 488540 18566 488592 18572
rect 488552 3482 488580 18566
rect 491312 3482 491340 120090
rect 487172 3454 488212 3482
rect 488552 3454 489408 3482
rect 491312 3454 491800 3482
rect 486974 3431 487030 3440
rect 486988 480 487016 3431
rect 488184 480 488212 3454
rect 489380 480 489408 3454
rect 490564 2848 490616 2854
rect 490564 2790 490616 2796
rect 490576 480 490604 2790
rect 491772 480 491800 3454
rect 492692 3346 492720 264182
rect 494072 3482 494100 266591
rect 511998 265432 512054 265441
rect 511998 265367 512054 265376
rect 498200 264104 498252 264110
rect 498200 264046 498252 264052
rect 497464 225004 497516 225010
rect 497464 224946 497516 224952
rect 496084 67652 496136 67658
rect 496084 67594 496136 67600
rect 494704 57996 494756 58002
rect 494704 57938 494756 57944
rect 494716 41410 494744 57938
rect 494704 41404 494756 41410
rect 494704 41346 494756 41352
rect 495348 6452 495400 6458
rect 495348 6394 495400 6400
rect 494072 3454 494192 3482
rect 492692 3318 492996 3346
rect 492968 480 492996 3318
rect 494164 480 494192 3454
rect 495360 480 495388 6394
rect 496096 3602 496124 67594
rect 496084 3596 496136 3602
rect 496084 3538 496136 3544
rect 497476 3466 497504 224946
rect 497740 3664 497792 3670
rect 497740 3606 497792 3612
rect 496544 3460 496596 3466
rect 496544 3402 496596 3408
rect 497464 3460 497516 3466
rect 497464 3402 497516 3408
rect 496556 480 496584 3402
rect 497752 480 497780 3606
rect 498212 3482 498240 264046
rect 499580 263152 499632 263158
rect 499580 263094 499632 263100
rect 499592 3482 499620 263094
rect 502984 176724 503036 176730
rect 502984 176666 503036 176672
rect 501604 164280 501656 164286
rect 501604 164222 501656 164228
rect 501616 88330 501644 164222
rect 501604 88324 501656 88330
rect 501604 88266 501656 88272
rect 502432 28280 502484 28286
rect 502432 28222 502484 28228
rect 500960 25628 501012 25634
rect 500960 25570 501012 25576
rect 500972 3482 501000 25570
rect 502444 3602 502472 28222
rect 502996 3738 503024 176666
rect 506480 44192 506532 44198
rect 506480 44134 506532 44140
rect 505100 17332 505152 17338
rect 505100 17274 505152 17280
rect 502984 3732 503036 3738
rect 502984 3674 503036 3680
rect 502340 3596 502392 3602
rect 502340 3538 502392 3544
rect 502432 3596 502484 3602
rect 502432 3538 502484 3544
rect 503628 3596 503680 3602
rect 503628 3538 503680 3544
rect 502352 3482 502380 3538
rect 498212 3454 498976 3482
rect 499592 3454 500172 3482
rect 500972 3454 501276 3482
rect 502352 3454 502472 3482
rect 498948 480 498976 3454
rect 500144 480 500172 3454
rect 501248 480 501276 3454
rect 502444 480 502472 3454
rect 503640 480 503668 3538
rect 505112 3482 505140 17274
rect 506492 3482 506520 44134
rect 510620 15904 510672 15910
rect 510620 15846 510672 15852
rect 507860 11824 507912 11830
rect 507860 11766 507912 11772
rect 507872 3482 507900 11766
rect 510632 3482 510660 15846
rect 505112 3454 506060 3482
rect 506492 3454 507256 3482
rect 507872 3454 508452 3482
rect 504822 3360 504878 3369
rect 504822 3295 504878 3304
rect 504836 480 504864 3295
rect 506032 480 506060 3454
rect 507228 480 507256 3454
rect 508424 480 508452 3454
rect 509608 3460 509660 3466
rect 510632 3454 510844 3482
rect 509608 3402 509660 3408
rect 509620 480 509648 3402
rect 510816 480 510844 3454
rect 512012 480 512040 265367
rect 514024 215348 514076 215354
rect 514024 215290 514076 215296
rect 512090 36544 512146 36553
rect 512090 36479 512146 36488
rect 512104 3482 512132 36479
rect 513380 17264 513432 17270
rect 513380 17206 513432 17212
rect 513392 3618 513420 17206
rect 514036 4146 514064 215290
rect 517520 193248 517572 193254
rect 517520 193190 517572 193196
rect 516140 19984 516192 19990
rect 516140 19926 516192 19932
rect 514760 18692 514812 18698
rect 514760 18634 514812 18640
rect 514024 4140 514076 4146
rect 514024 4082 514076 4088
rect 514576 4140 514628 4146
rect 514576 4082 514628 4088
rect 513392 3590 514432 3618
rect 512104 3454 513236 3482
rect 513208 480 513236 3454
rect 514404 480 514432 3590
rect 514588 3466 514616 4082
rect 514772 3482 514800 18634
rect 516152 3482 516180 19926
rect 517532 3482 517560 193190
rect 518912 3482 518940 267990
rect 520292 3670 520320 269894
rect 521660 267844 521712 267850
rect 521660 267786 521712 267792
rect 520372 18760 520424 18766
rect 520372 18702 520424 18708
rect 520280 3664 520332 3670
rect 520280 3606 520332 3612
rect 520384 3482 520412 18702
rect 521476 3664 521528 3670
rect 521476 3606 521528 3612
rect 514576 3460 514628 3466
rect 514772 3454 515628 3482
rect 516152 3454 516824 3482
rect 517532 3454 517928 3482
rect 518912 3454 519124 3482
rect 514576 3402 514628 3408
rect 515600 480 515628 3454
rect 516796 480 516824 3454
rect 517900 480 517928 3454
rect 519096 480 519124 3454
rect 520292 3454 520412 3482
rect 520292 480 520320 3454
rect 521488 480 521516 3606
rect 521672 3482 521700 267786
rect 528558 265296 528614 265305
rect 528558 265231 528614 265240
rect 527180 263628 527232 263634
rect 527180 263570 527232 263576
rect 526258 6760 526314 6769
rect 526258 6695 526314 6704
rect 523868 4956 523920 4962
rect 523868 4898 523920 4904
rect 521672 3454 522712 3482
rect 522684 480 522712 3454
rect 523880 480 523908 4898
rect 525062 4856 525118 4865
rect 525062 4791 525118 4800
rect 525076 480 525104 4791
rect 526272 480 526300 6695
rect 527192 3482 527220 263570
rect 528572 3482 528600 265231
rect 531318 264208 531374 264217
rect 531318 264143 531374 264152
rect 529938 32600 529994 32609
rect 529938 32535 529994 32544
rect 528652 16108 528704 16114
rect 528652 16050 528704 16056
rect 528664 3670 528692 16050
rect 528652 3664 528704 3670
rect 528652 3606 528704 3612
rect 529848 3664 529900 3670
rect 529848 3606 529900 3612
rect 527192 3454 527496 3482
rect 528572 3454 528692 3482
rect 527468 480 527496 3454
rect 528664 480 528692 3454
rect 529860 480 529888 3606
rect 529952 3482 529980 32535
rect 531332 3482 531360 264143
rect 533356 40050 533384 700266
rect 543568 698290 543596 703446
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 542728 698284 542780 698290
rect 542728 698226 542780 698232
rect 543556 698284 543608 698290
rect 543556 698226 543608 698232
rect 542740 688702 542768 698226
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 542728 688696 542780 688702
rect 542728 688638 542780 688644
rect 542544 688628 542596 688634
rect 542544 688570 542596 688576
rect 542556 685930 542584 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 542464 685902 542584 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 542464 684486 542492 685902
rect 580172 685850 580224 685856
rect 542452 684480 542504 684486
rect 542452 684422 542504 684428
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 542820 666596 542872 666602
rect 542820 666538 542872 666544
rect 542832 659682 542860 666538
rect 542648 659654 542860 659682
rect 542648 647290 542676 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 542544 647284 542596 647290
rect 542544 647226 542596 647232
rect 542636 647284 542688 647290
rect 542636 647226 542688 647232
rect 542556 640422 542584 647226
rect 542544 640416 542596 640422
rect 542544 640358 542596 640364
rect 542636 640416 542688 640422
rect 542636 640358 542688 640364
rect 542648 630698 542676 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 542452 630692 542504 630698
rect 542452 630634 542504 630640
rect 542636 630692 542688 630698
rect 542636 630634 542688 630640
rect 542464 630578 542492 630634
rect 542464 630550 542584 630578
rect 542556 621058 542584 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 542556 621030 542676 621058
rect 542648 611386 542676 621030
rect 542452 611380 542504 611386
rect 542452 611322 542504 611328
rect 542636 611380 542688 611386
rect 542636 611322 542688 611328
rect 542464 611266 542492 611322
rect 542464 611238 542584 611266
rect 542556 608598 542584 611238
rect 542544 608592 542596 608598
rect 542544 608534 542596 608540
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 542728 601724 542780 601730
rect 542728 601666 542780 601672
rect 542740 598942 542768 601666
rect 542728 598936 542780 598942
rect 542728 598878 542780 598884
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 542820 589348 542872 589354
rect 542820 589290 542872 589296
rect 542832 582486 542860 589290
rect 542820 582480 542872 582486
rect 542820 582422 542872 582428
rect 542728 582344 542780 582350
rect 542728 582286 542780 582292
rect 542740 572642 542768 582286
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 542556 572614 542768 572642
rect 542556 569922 542584 572614
rect 542464 569894 542584 569922
rect 542464 563174 542492 569894
rect 542452 563168 542504 563174
rect 542452 563110 542504 563116
rect 542452 563032 542504 563038
rect 542452 562974 542504 562980
rect 542464 560250 542492 562974
rect 542452 560244 542504 560250
rect 542452 560186 542504 560192
rect 534078 556608 534134 556617
rect 534078 556543 534134 556552
rect 540978 556608 541034 556617
rect 540978 556543 541034 556552
rect 533986 556200 534042 556209
rect 534092 556186 534120 556543
rect 540992 556209 541020 556543
rect 553398 556472 553454 556481
rect 553320 556430 553398 556458
rect 553320 556345 553348 556430
rect 553398 556407 553454 556416
rect 553306 556336 553362 556345
rect 553306 556271 553362 556280
rect 534042 556158 534120 556186
rect 540978 556200 541034 556209
rect 533986 556135 534042 556144
rect 540978 556135 541034 556144
rect 542636 550656 542688 550662
rect 542636 550598 542688 550604
rect 542648 543658 542676 550598
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 542452 543652 542504 543658
rect 542452 543594 542504 543600
rect 542636 543652 542688 543658
rect 542636 543594 542688 543600
rect 542464 534070 542492 543594
rect 542452 534064 542504 534070
rect 542452 534006 542504 534012
rect 542636 534064 542688 534070
rect 542636 534006 542688 534012
rect 542648 524482 542676 534006
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 542636 524476 542688 524482
rect 542636 524418 542688 524424
rect 542728 524408 542780 524414
rect 542728 524350 542780 524356
rect 542740 521665 542768 524350
rect 542542 521656 542598 521665
rect 542542 521591 542598 521600
rect 542726 521656 542782 521665
rect 542726 521591 542782 521600
rect 542556 512038 542584 521591
rect 542544 512032 542596 512038
rect 542544 511974 542596 511980
rect 542820 512032 542872 512038
rect 542820 511974 542872 511980
rect 542832 502382 542860 511974
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 542636 502376 542688 502382
rect 542358 502344 542414 502353
rect 542358 502279 542414 502288
rect 542634 502344 542636 502353
rect 542820 502376 542872 502382
rect 542688 502344 542690 502353
rect 542820 502318 542872 502324
rect 542634 502279 542690 502288
rect 542372 492697 542400 502279
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 542358 492688 542414 492697
rect 542358 492623 542414 492632
rect 542542 492688 542598 492697
rect 542542 492623 542544 492632
rect 542596 492623 542598 492632
rect 542544 492594 542596 492600
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 542544 485784 542596 485790
rect 542544 485726 542596 485732
rect 542556 483018 542584 485726
rect 542556 482990 542676 483018
rect 542648 476134 542676 482990
rect 542452 476128 542504 476134
rect 542636 476128 542688 476134
rect 542504 476076 542584 476082
rect 542452 476070 542584 476076
rect 542636 476070 542688 476076
rect 542464 476054 542584 476070
rect 542556 473346 542584 476054
rect 542544 473340 542596 473346
rect 542544 473282 542596 473288
rect 542544 466404 542596 466410
rect 542544 466346 542596 466352
rect 542556 463706 542584 466346
rect 542556 463678 542676 463706
rect 542648 454073 542676 463678
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 542358 454064 542414 454073
rect 542358 453999 542414 454008
rect 542634 454064 542690 454073
rect 542634 453999 542690 454008
rect 542372 447166 542400 453999
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580184 451314 580212 451687
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 542360 447160 542412 447166
rect 542360 447102 542412 447108
rect 542452 447092 542504 447098
rect 542452 447034 542504 447040
rect 542464 444378 542492 447034
rect 542176 444372 542228 444378
rect 542176 444314 542228 444320
rect 542452 444372 542504 444378
rect 542452 444314 542504 444320
rect 542188 434761 542216 444314
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 542174 434752 542230 434761
rect 542174 434687 542230 434696
rect 542358 434752 542414 434761
rect 542358 434687 542414 434696
rect 542372 427854 542400 434687
rect 542360 427848 542412 427854
rect 542360 427790 542412 427796
rect 542452 427780 542504 427786
rect 542452 427722 542504 427728
rect 542464 425066 542492 427722
rect 542176 425060 542228 425066
rect 542176 425002 542228 425008
rect 542452 425060 542504 425066
rect 542452 425002 542504 425008
rect 542188 415449 542216 425002
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 580184 415478 580212 416463
rect 580172 415472 580224 415478
rect 542174 415440 542230 415449
rect 542174 415375 542230 415384
rect 542358 415440 542414 415449
rect 580172 415414 580224 415420
rect 542358 415375 542414 415384
rect 542372 408542 542400 415375
rect 542360 408536 542412 408542
rect 542360 408478 542412 408484
rect 542452 408400 542504 408406
rect 542452 408342 542504 408348
rect 542464 405686 542492 408342
rect 542452 405680 542504 405686
rect 542452 405622 542504 405628
rect 580170 404832 580226 404841
rect 580170 404767 580226 404776
rect 580184 404394 580212 404767
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 542452 398812 542504 398818
rect 542452 398754 542504 398760
rect 542464 389230 542492 398754
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 580184 392018 580212 392935
rect 580172 392012 580224 392018
rect 580172 391954 580224 391960
rect 542452 389224 542504 389230
rect 542452 389166 542504 389172
rect 542452 389088 542504 389094
rect 542452 389030 542504 389036
rect 542464 379506 542492 389030
rect 542452 379500 542504 379506
rect 542452 379442 542504 379448
rect 542636 379500 542688 379506
rect 542636 379442 542688 379448
rect 542648 371906 542676 379442
rect 542648 371878 542768 371906
rect 542740 357542 542768 371878
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580184 368558 580212 369543
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 580170 357912 580226 357921
rect 580170 357847 580226 357856
rect 542728 357536 542780 357542
rect 542728 357478 542780 357484
rect 580184 357474 580212 357847
rect 580172 357468 580224 357474
rect 580172 357410 580224 357416
rect 542728 353388 542780 353394
rect 542728 353330 542780 353336
rect 542740 353274 542768 353330
rect 542740 353258 542860 353274
rect 542740 353252 542872 353258
rect 542740 353246 542820 353252
rect 542820 353194 542872 353200
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580184 345098 580212 346015
rect 580172 345092 580224 345098
rect 580172 345034 580224 345040
rect 542820 340808 542872 340814
rect 542820 340750 542872 340756
rect 542832 331514 542860 340750
rect 542740 331486 542860 331514
rect 542740 325718 542768 331486
rect 542636 325712 542688 325718
rect 542636 325654 542688 325660
rect 542728 325712 542780 325718
rect 542728 325654 542780 325660
rect 542648 318850 542676 325654
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 580184 321638 580212 322623
rect 580172 321632 580224 321638
rect 580172 321574 580224 321580
rect 542544 318844 542596 318850
rect 542544 318786 542596 318792
rect 542636 318844 542688 318850
rect 542636 318786 542688 318792
rect 542556 311982 542584 318786
rect 542544 311976 542596 311982
rect 542544 311918 542596 311924
rect 542636 311976 542688 311982
rect 542636 311918 542688 311924
rect 542648 302258 542676 311918
rect 579802 310856 579858 310865
rect 579802 310791 579858 310800
rect 579816 310554 579844 310791
rect 579804 310548 579856 310554
rect 579804 310490 579856 310496
rect 542452 302252 542504 302258
rect 542452 302194 542504 302200
rect 542636 302252 542688 302258
rect 542636 302194 542688 302200
rect 542464 302138 542492 302194
rect 542464 302110 542584 302138
rect 542556 292618 542584 302110
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 580184 298178 580212 299095
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 542556 292590 542676 292618
rect 542648 289814 542676 292590
rect 542636 289808 542688 289814
rect 542636 289750 542688 289756
rect 542452 280220 542504 280226
rect 542452 280162 542504 280168
rect 542464 273306 542492 280162
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580184 274718 580212 275703
rect 580172 274712 580224 274718
rect 580172 274654 580224 274660
rect 542464 273278 542676 273306
rect 542452 268660 542504 268666
rect 542452 268602 542504 268608
rect 539600 267912 539652 267918
rect 539600 267854 539652 267860
rect 535460 244316 535512 244322
rect 535460 244258 535512 244264
rect 534080 43512 534132 43518
rect 534080 43454 534132 43460
rect 533344 40044 533396 40050
rect 533344 39986 533396 39992
rect 532700 17468 532752 17474
rect 532700 17410 532752 17416
rect 532712 3482 532740 17410
rect 534092 3482 534120 43454
rect 535472 3482 535500 244258
rect 538220 51740 538272 51746
rect 538220 51682 538272 51688
rect 538128 7744 538180 7750
rect 538128 7686 538180 7692
rect 536930 3496 536986 3505
rect 529952 3454 531084 3482
rect 531332 3454 532280 3482
rect 532712 3454 533476 3482
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 531056 480 531084 3454
rect 532252 480 532280 3454
rect 533448 480 533476 3454
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536930 3431 536986 3440
rect 536944 480 536972 3431
rect 538140 480 538168 7686
rect 538232 3482 538260 51682
rect 539612 3482 539640 267854
rect 542360 267776 542412 267782
rect 542360 267718 542412 267724
rect 542372 244254 542400 267718
rect 542360 244248 542412 244254
rect 542360 244190 542412 244196
rect 542358 231840 542414 231849
rect 542358 231775 542414 231784
rect 542372 222222 542400 231775
rect 542360 222216 542412 222222
rect 542360 222158 542412 222164
rect 542360 169108 542412 169114
rect 542360 169050 542412 169056
rect 542372 161430 542400 169050
rect 542360 161424 542412 161430
rect 542360 161366 542412 161372
rect 542360 151836 542412 151842
rect 542360 151778 542412 151784
rect 542372 142118 542400 151778
rect 542360 142112 542412 142118
rect 542360 142054 542412 142060
rect 542360 132524 542412 132530
rect 542360 132466 542412 132472
rect 542372 128314 542400 132466
rect 542360 128308 542412 128314
rect 542360 128250 542412 128256
rect 542360 115932 542412 115938
rect 542360 115874 542412 115880
rect 542372 106321 542400 115874
rect 542358 106312 542414 106321
rect 542358 106247 542414 106256
rect 541716 6248 541768 6254
rect 541716 6190 541768 6196
rect 538232 3454 539364 3482
rect 539612 3454 540560 3482
rect 539336 480 539364 3454
rect 540532 480 540560 3454
rect 541728 480 541756 6190
rect 542464 3482 542492 268602
rect 542648 267782 542676 273278
rect 579804 267980 579856 267986
rect 579804 267922 579856 267928
rect 542636 267776 542688 267782
rect 542636 267718 542688 267724
rect 554778 265840 554834 265849
rect 554778 265775 554834 265784
rect 547880 265056 547932 265062
rect 547880 264998 547932 265004
rect 543738 264480 543794 264489
rect 543738 264415 543794 264424
rect 542636 244248 542688 244254
rect 542636 244190 542688 244196
rect 542648 234682 542676 244190
rect 542648 234654 542768 234682
rect 542740 231878 542768 234654
rect 542544 231872 542596 231878
rect 542542 231840 542544 231849
rect 542728 231872 542780 231878
rect 542596 231840 542598 231849
rect 542728 231814 542780 231820
rect 542542 231775 542598 231784
rect 542636 222216 542688 222222
rect 542636 222158 542688 222164
rect 542648 215370 542676 222158
rect 542648 215342 542768 215370
rect 542740 212537 542768 215342
rect 542542 212528 542598 212537
rect 542542 212463 542598 212472
rect 542726 212528 542782 212537
rect 542726 212463 542782 212472
rect 542556 202910 542584 212463
rect 542544 202904 542596 202910
rect 542544 202846 542596 202852
rect 542636 202904 542688 202910
rect 542636 202846 542688 202852
rect 542648 196042 542676 202846
rect 542636 196036 542688 196042
rect 542636 195978 542688 195984
rect 542728 195968 542780 195974
rect 542728 195910 542780 195916
rect 542740 193225 542768 195910
rect 542542 193216 542598 193225
rect 542542 193151 542598 193160
rect 542726 193216 542782 193225
rect 542726 193151 542782 193160
rect 542556 183598 542584 193151
rect 542544 183592 542596 183598
rect 542544 183534 542596 183540
rect 542820 183592 542872 183598
rect 542820 183534 542872 183540
rect 542832 173942 542860 183534
rect 542636 173936 542688 173942
rect 542636 173878 542688 173884
rect 542820 173936 542872 173942
rect 542820 173878 542872 173884
rect 542648 169114 542676 173878
rect 542636 169108 542688 169114
rect 542636 169050 542688 169056
rect 542636 161424 542688 161430
rect 542636 161366 542688 161372
rect 542648 151842 542676 161366
rect 542636 151836 542688 151842
rect 542636 151778 542688 151784
rect 542636 142112 542688 142118
rect 542636 142054 542688 142060
rect 542648 132530 542676 142054
rect 542636 132524 542688 132530
rect 542636 132466 542688 132472
rect 542636 128308 542688 128314
rect 542636 128250 542688 128256
rect 542648 120714 542676 128250
rect 542648 120686 542768 120714
rect 542740 115977 542768 120686
rect 542542 115968 542598 115977
rect 542542 115903 542544 115912
rect 542596 115903 542598 115912
rect 542726 115968 542782 115977
rect 542726 115903 542782 115912
rect 542544 115874 542596 115880
rect 542634 106312 542690 106321
rect 542634 106247 542690 106256
rect 542648 101454 542676 106247
rect 542636 101448 542688 101454
rect 542636 101390 542688 101396
rect 542728 99340 542780 99346
rect 542728 99282 542780 99288
rect 542740 89706 542768 99282
rect 542648 89678 542768 89706
rect 542648 80073 542676 89678
rect 542634 80064 542690 80073
rect 542634 79999 542690 80008
rect 542634 77344 542690 77353
rect 542634 77279 542690 77288
rect 542648 77217 542676 77279
rect 542634 77208 542690 77217
rect 542634 77143 542690 77152
rect 542542 67688 542598 67697
rect 542542 67623 542598 67632
rect 542556 67590 542584 67623
rect 542544 67584 542596 67590
rect 542544 67526 542596 67532
rect 542728 67584 542780 67590
rect 542728 67526 542780 67532
rect 542740 60602 542768 67526
rect 542648 60574 542768 60602
rect 542648 42129 542676 60574
rect 542634 42120 542690 42129
rect 542634 42055 542690 42064
rect 543752 3482 543780 264415
rect 546500 31136 546552 31142
rect 546500 31078 546552 31084
rect 545304 7812 545356 7818
rect 545304 7754 545356 7760
rect 542464 3454 542952 3482
rect 543752 3454 544148 3482
rect 542924 480 542952 3454
rect 544120 480 544148 3454
rect 545316 480 545344 7754
rect 546512 480 546540 31078
rect 546592 21412 546644 21418
rect 546592 21354 546644 21360
rect 546604 3482 546632 21354
rect 546604 3454 547736 3482
rect 547708 480 547736 3454
rect 547892 610 547920 264998
rect 554044 99408 554096 99414
rect 554044 99350 554096 99356
rect 549258 15872 549314 15881
rect 549258 15807 549314 15816
rect 549272 610 549300 15807
rect 554056 13122 554084 99350
rect 553400 13116 553452 13122
rect 553400 13058 553452 13064
rect 554044 13116 554096 13122
rect 554044 13058 554096 13064
rect 551192 5024 551244 5030
rect 551192 4966 551244 4972
rect 547880 604 547932 610
rect 547880 546 547932 552
rect 548892 604 548944 610
rect 548892 546 548944 552
rect 549260 604 549312 610
rect 549260 546 549312 552
rect 550088 604 550140 610
rect 550088 546 550140 552
rect 548904 480 548932 546
rect 550100 480 550128 546
rect 551204 480 551232 4966
rect 552388 3596 552440 3602
rect 552388 3538 552440 3544
rect 552400 480 552428 3538
rect 553412 626 553440 13058
rect 553412 598 553624 626
rect 553596 480 553624 598
rect 554792 480 554820 265775
rect 565818 265568 565874 265577
rect 565818 265503 565874 265512
rect 556160 263220 556212 263226
rect 556160 263162 556212 263168
rect 555976 7608 556028 7614
rect 555976 7550 556028 7556
rect 555988 480 556016 7550
rect 556172 610 556200 263162
rect 561680 47592 561732 47598
rect 561680 47534 561732 47540
rect 558920 26920 558972 26926
rect 558920 26862 558972 26868
rect 558366 6624 558422 6633
rect 558366 6559 558422 6568
rect 556160 604 556212 610
rect 556160 546 556212 552
rect 557172 604 557224 610
rect 557172 546 557224 552
rect 557184 480 557212 546
rect 558380 480 558408 6559
rect 558932 3482 558960 26862
rect 560300 13116 560352 13122
rect 560300 13058 560352 13064
rect 560312 3482 560340 13058
rect 561692 3482 561720 47534
rect 563060 29640 563112 29646
rect 563060 29582 563112 29588
rect 563072 3482 563100 29582
rect 563150 24168 563206 24177
rect 563150 24103 563206 24112
rect 563164 3602 563192 24103
rect 565542 6488 565598 6497
rect 565542 6423 565598 6432
rect 563152 3596 563204 3602
rect 563152 3538 563204 3544
rect 564348 3596 564400 3602
rect 564348 3538 564400 3544
rect 558932 3454 559604 3482
rect 560312 3454 560800 3482
rect 561692 3454 561996 3482
rect 563072 3454 563192 3482
rect 559576 480 559604 3454
rect 560772 480 560800 3454
rect 561968 480 561996 3454
rect 563164 480 563192 3454
rect 564360 480 564388 3538
rect 565556 480 565584 6423
rect 565832 3482 565860 265503
rect 574742 265160 574798 265169
rect 574742 265095 574798 265104
rect 572720 33788 572772 33794
rect 572720 33730 572772 33736
rect 571338 32464 571394 32473
rect 571338 32399 571394 32408
rect 569960 14476 570012 14482
rect 569960 14418 570012 14424
rect 569038 6352 569094 6361
rect 569038 6287 569094 6296
rect 567844 3528 567896 3534
rect 565832 3454 566780 3482
rect 567844 3470 567896 3476
rect 566752 480 566780 3454
rect 567856 480 567884 3470
rect 569052 480 569080 6287
rect 569972 3482 570000 14418
rect 571352 3482 571380 32399
rect 572626 6216 572682 6225
rect 572626 6151 572682 6160
rect 569972 3454 570276 3482
rect 571352 3454 571472 3482
rect 570248 480 570276 3454
rect 571444 480 571472 3454
rect 572640 480 572668 6151
rect 572732 3482 572760 33730
rect 574756 3534 574784 265095
rect 579816 263945 579844 267922
rect 581090 264344 581146 264353
rect 581090 264279 581146 264288
rect 579802 263936 579858 263945
rect 579802 263871 579858 263880
rect 575478 263800 575534 263809
rect 575478 263735 575534 263744
rect 575020 8968 575072 8974
rect 575020 8910 575072 8916
rect 574744 3528 574796 3534
rect 572732 3454 573864 3482
rect 574744 3470 574796 3476
rect 573836 480 573864 3454
rect 575032 480 575060 8910
rect 575492 3482 575520 263735
rect 578240 253224 578292 253230
rect 578240 253166 578292 253172
rect 575492 3454 576256 3482
rect 576228 480 576256 3454
rect 577412 3460 577464 3466
rect 577412 3402 577464 3408
rect 577424 480 577452 3402
rect 578252 626 578280 253166
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 580262 228848 580318 228857
rect 580262 228783 580318 228792
rect 579894 205320 579950 205329
rect 579894 205255 579950 205264
rect 579908 204338 579936 205255
rect 579896 204332 579948 204338
rect 579896 204274 579948 204280
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 580184 169794 580212 170031
rect 580172 169788 580224 169794
rect 580172 169730 580224 169736
rect 579894 158400 579950 158409
rect 579894 158335 579950 158344
rect 579908 157418 579936 158335
rect 579896 157412 579948 157418
rect 579896 157354 579948 157360
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580184 133958 580212 134807
rect 580172 133952 580224 133958
rect 580172 133894 580224 133900
rect 579896 124160 579948 124166
rect 579896 124102 579948 124108
rect 579908 123185 579936 124102
rect 579894 123176 579950 123185
rect 579894 123111 579950 123120
rect 579896 88324 579948 88330
rect 579896 88266 579948 88272
rect 579908 87961 579936 88266
rect 579894 87952 579950 87961
rect 579894 87887 579950 87896
rect 579620 77240 579672 77246
rect 579620 77182 579672 77188
rect 579632 76265 579660 77182
rect 579618 76256 579674 76265
rect 579618 76191 579674 76200
rect 580172 64864 580224 64870
rect 580172 64806 580224 64812
rect 580184 64569 580212 64806
rect 580170 64560 580226 64569
rect 580170 64495 580226 64504
rect 580276 42090 580304 228783
rect 580264 42084 580316 42090
rect 580264 42026 580316 42032
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 579804 4820 579856 4826
rect 579804 4762 579856 4768
rect 578252 598 578648 626
rect 578620 480 578648 598
rect 579816 480 579844 4762
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581012 480 581040 3470
rect 581104 610 581132 264279
rect 581092 604 581144 610
rect 581092 546 581144 552
rect 582196 604 582248 610
rect 582196 546 582248 552
rect 582208 480 582236 546
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3330 682216 3386 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3330 653520 3386 653576
rect 3330 652840 3386 652896
rect 4066 624824 4122 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 4066 567296 4122 567352
rect 4066 553016 4122 553072
rect 3974 538600 4030 538656
rect 3882 509904 3938 509960
rect 4066 495508 4122 495544
rect 4066 495488 4068 495508
rect 4068 495488 4120 495508
rect 4120 495488 4122 495508
rect 3330 481072 3386 481128
rect 3422 452376 3478 452432
rect 3146 294344 3202 294400
rect 2962 222536 3018 222592
rect 3330 165008 3386 165064
rect 2778 122032 2834 122088
rect 3790 437960 3846 438016
rect 4066 423700 4122 423736
rect 4066 423680 4068 423700
rect 4068 423680 4120 423700
rect 4120 423680 4122 423700
rect 4066 394984 4122 395040
rect 3974 380568 4030 380624
rect 4066 366152 4122 366208
rect 4066 337456 4122 337512
rect 3606 323040 3662 323096
rect 4066 308760 4122 308816
rect 3698 280064 3754 280120
rect 3882 265648 3938 265704
rect 4066 251252 4122 251288
rect 4066 251232 4068 251252
rect 4068 251232 4120 251252
rect 4120 251232 4122 251252
rect 4066 236952 4122 237008
rect 4066 180648 4122 180704
rect 4066 179424 4122 179480
rect 3606 150728 3662 150784
rect 3514 64504 3570 64560
rect 3514 50088 3570 50144
rect 3974 136312 4030 136368
rect 4066 107652 4068 107672
rect 4068 107652 4120 107672
rect 4120 107652 4122 107672
rect 4066 107616 4122 107652
rect 3974 78920 4030 78976
rect 8114 531256 8170 531312
rect 8390 531256 8446 531312
rect 8114 511944 8170 512000
rect 8390 511944 8446 512000
rect 7930 482976 7986 483032
rect 8206 482976 8262 483032
rect 7838 434696 7894 434752
rect 8022 434696 8078 434752
rect 4894 194520 4950 194576
rect 4894 193840 4950 193896
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3146 21392 3202 21448
rect 12346 194520 12402 194576
rect 12530 194384 12586 194440
rect 22190 194520 22246 194576
rect 27618 194540 27674 194576
rect 27618 194520 27620 194540
rect 27620 194520 27672 194540
rect 27672 194520 27674 194540
rect 22006 194384 22062 194440
rect 37186 194248 37242 194304
rect 53470 8880 53526 8936
rect 2962 7112 3018 7168
rect 54758 9016 54814 9072
rect 55862 6704 55918 6760
rect 56046 6296 56102 6352
rect 56138 3984 56194 4040
rect 57334 142024 57390 142080
rect 57242 6160 57298 6216
rect 57334 3440 57390 3496
rect 59358 260344 59414 260400
rect 59266 239944 59322 240000
rect 59174 233960 59230 234016
rect 59082 229608 59138 229664
rect 58898 187176 58954 187232
rect 58806 174120 58862 174176
rect 58714 146376 58770 146432
rect 58622 119992 58678 120048
rect 58990 185816 59046 185872
rect 59358 222264 59414 222320
rect 59358 220904 59414 220960
rect 59450 217912 59506 217968
rect 59358 216588 59360 216608
rect 59360 216588 59412 216608
rect 59412 216588 59414 216608
rect 59358 216552 59414 216588
rect 59358 214920 59414 214976
rect 59358 213560 59414 213616
rect 59358 206216 59414 206272
rect 59358 203224 59414 203280
rect 59358 198872 59414 198928
rect 59358 194520 59414 194576
rect 60462 257352 60518 257408
rect 60462 236952 60518 237008
rect 60370 193160 60426 193216
rect 60278 190168 60334 190224
rect 59358 188808 59414 188864
rect 59910 182824 59966 182880
rect 59358 181464 59414 181520
rect 59542 175480 59598 175536
rect 59358 168136 59414 168192
rect 59358 165416 59414 165472
rect 60094 153720 60150 153776
rect 59358 150728 59414 150784
rect 59358 143384 59414 143440
rect 59358 131688 59414 131744
rect 59726 130328 59782 130384
rect 59358 128696 59414 128752
rect 59358 121352 59414 121408
rect 59358 118632 59414 118688
rect 59634 112648 59690 112704
rect 59358 103944 59414 104000
rect 59358 100952 59414 101008
rect 60186 133048 60242 133104
rect 59358 90888 59414 90944
rect 59726 87896 59782 87952
rect 59634 83544 59690 83600
rect 59358 77560 59414 77616
rect 59358 74588 59414 74624
rect 59358 74568 59360 74588
rect 59360 74568 59412 74588
rect 59412 74568 59414 74588
rect 59358 65864 59414 65920
rect 59358 60152 59414 60208
rect 60278 122984 60334 123040
rect 60278 105304 60334 105360
rect 60186 81504 60242 81560
rect 60002 80552 60058 80608
rect 59910 64504 59966 64560
rect 60094 79192 60150 79248
rect 60738 253000 60794 253056
rect 60646 172760 60702 172816
rect 60554 149368 60610 149424
rect 60646 111288 60702 111344
rect 60646 106936 60702 106992
rect 60554 97688 60610 97744
rect 60462 75792 60518 75848
rect 60462 49544 60518 49600
rect 60830 250008 60886 250064
rect 61014 251640 61070 251696
rect 60922 238312 60978 238368
rect 60922 219544 60978 219600
rect 61106 248648 61162 248704
rect 61106 208256 61162 208312
rect 61106 163784 61162 163840
rect 61014 73072 61070 73128
rect 61014 70216 61070 70272
rect 61290 223896 61346 223952
rect 62394 205808 62450 205864
rect 62394 201456 62450 201512
rect 61290 193296 61346 193352
rect 61290 191528 61346 191584
rect 61198 159432 61254 159488
rect 61198 94696 61254 94752
rect 64970 265376 65026 265432
rect 74906 269184 74962 269240
rect 86682 268368 86738 268424
rect 78770 267144 78826 267200
rect 79874 265240 79930 265296
rect 88706 265784 88762 265840
rect 102506 267824 102562 267880
rect 103610 266736 103666 266792
rect 107474 266872 107530 266928
rect 106554 266464 106610 266520
rect 114466 265104 114522 265160
rect 126978 265512 127034 265568
rect 129186 266464 129242 266520
rect 142066 266600 142122 266656
rect 149058 266872 149114 266928
rect 63222 264288 63278 264344
rect 113546 264288 113602 264344
rect 170310 700440 170366 700496
rect 218978 700304 219034 700360
rect 199474 269320 199530 269376
rect 200394 267960 200450 268016
rect 246026 269592 246082 269648
rect 244922 269456 244978 269512
rect 209686 264424 209742 264480
rect 238114 267008 238170 267064
rect 241058 265648 241114 265704
rect 267646 700304 267702 700360
rect 257802 266328 257858 266384
rect 159546 264288 159602 264344
rect 163410 264288 163466 264344
rect 201682 264288 201738 264344
rect 222566 264288 222622 264344
rect 264794 267280 264850 267336
rect 263598 266600 263654 266656
rect 270498 266600 270554 266656
rect 271786 266328 271842 266384
rect 271786 264968 271842 265024
rect 281078 267008 281134 267064
rect 268290 264560 268346 264616
rect 279882 264560 279938 264616
rect 255134 264288 255190 264344
rect 259458 264288 259514 264344
rect 268290 264288 268346 264344
rect 275006 264288 275062 264344
rect 279882 264288 279938 264344
rect 280986 263472 281042 263528
rect 280986 172488 281042 172544
rect 280986 154536 281042 154592
rect 62394 128152 62450 128208
rect 280986 135244 281042 135280
rect 280986 135224 280988 135244
rect 280988 135224 281040 135244
rect 281040 135224 281042 135244
rect 62394 116048 62450 116104
rect 62394 111424 62450 111480
rect 62394 106256 62450 106312
rect 62210 105984 62266 106040
rect 62210 98232 62266 98288
rect 61382 97960 61438 98016
rect 61382 97688 61438 97744
rect 62394 93744 62450 93800
rect 62394 88576 62450 88632
rect 61382 86264 61438 86320
rect 281262 266736 281318 266792
rect 281170 219272 281226 219328
rect 281170 189624 281226 189680
rect 281354 154536 281410 154592
rect 281262 138488 281318 138544
rect 62394 81504 62450 81560
rect 62302 79872 62358 79928
rect 62210 70488 62266 70544
rect 62302 67768 62358 67824
rect 62210 60696 62266 60752
rect 61474 58520 61530 58576
rect 62026 46280 62082 46336
rect 62302 53896 62358 53952
rect 62210 44920 62266 44976
rect 281170 84360 281226 84416
rect 281078 60832 281134 60888
rect 281078 59608 281134 59664
rect 277030 43868 277032 43888
rect 277032 43868 277084 43888
rect 277084 43868 277086 43888
rect 277030 43832 277086 43868
rect 142066 43424 142122 43480
rect 79322 42744 79378 42800
rect 86314 42608 86370 42664
rect 96066 40840 96122 40896
rect 100114 41248 100170 41304
rect 101034 41112 101090 41168
rect 57426 3304 57482 3360
rect 121458 42064 121514 42120
rect 126610 3848 126666 3904
rect 136546 39208 136602 39264
rect 139306 29824 139362 29880
rect 146298 28192 146354 28248
rect 139674 3168 139730 3224
rect 150622 29008 150678 29064
rect 150806 29008 150862 29064
rect 153106 42200 153162 42256
rect 158442 42472 158498 42528
rect 161386 42336 161442 42392
rect 160006 15952 160062 16008
rect 168378 41112 168434 41168
rect 172978 6840 173034 6896
rect 171782 3712 171838 3768
rect 183558 30912 183614 30968
rect 190090 41928 190146 41984
rect 194506 39344 194562 39400
rect 200394 3576 200450 3632
rect 205914 42472 205970 42528
rect 209870 6024 209926 6080
rect 221738 40976 221794 41032
rect 232502 3576 232558 3632
rect 280066 3984 280122 4040
rect 281354 135360 281410 135416
rect 281630 129240 281686 129296
rect 281538 124888 281594 124944
rect 281630 104896 281686 104952
rect 281538 65320 281594 65376
rect 281998 185816 282054 185872
rect 281906 83544 281962 83600
rect 281906 62872 281962 62928
rect 282090 76200 282146 76256
rect 282366 92248 282422 92304
rect 282274 51176 282330 51232
rect 282918 235592 282974 235648
rect 282826 52400 282882 52456
rect 283194 261704 283250 261760
rect 283102 253000 283158 253056
rect 283010 209616 283066 209672
rect 283010 193160 283066 193216
rect 283194 241304 283250 241360
rect 283286 179832 283342 179888
rect 284114 251640 284170 251696
rect 284206 250008 284262 250064
rect 284206 248648 284262 248704
rect 284206 245676 284262 245712
rect 284206 245656 284208 245676
rect 284208 245656 284260 245676
rect 284260 245656 284262 245676
rect 284206 244316 284262 244352
rect 284206 244296 284208 244316
rect 284208 244296 284260 244316
rect 284260 244296 284262 244316
rect 283562 241440 283618 241496
rect 283838 238312 283894 238368
rect 283838 234776 283894 234832
rect 284206 233960 284262 234016
rect 283838 232056 283894 232112
rect 283562 231920 283618 231976
rect 284114 228248 284170 228304
rect 284206 226616 284262 226672
rect 284206 225256 284262 225312
rect 284206 217912 284262 217968
rect 284206 216552 284262 216608
rect 284206 213560 284262 213616
rect 284206 212200 284262 212256
rect 284114 207848 284170 207904
rect 284206 204856 284262 204912
rect 284206 201864 284262 201920
rect 284206 198872 284262 198928
rect 283562 197512 283618 197568
rect 283470 191528 283526 191584
rect 283378 161064 283434 161120
rect 283286 156440 283342 156496
rect 283378 152088 283434 152144
rect 284206 194520 284262 194576
rect 283838 192480 283894 192536
rect 284206 188808 284262 188864
rect 283930 184456 283986 184512
rect 283838 180376 283894 180432
rect 283838 165416 283894 165472
rect 283838 163784 283894 163840
rect 283838 149368 283894 149424
rect 283838 144744 283894 144800
rect 283838 143384 283894 143440
rect 283746 137672 283802 137728
rect 283470 127336 283526 127392
rect 283378 126928 283434 126984
rect 283378 125976 283434 126032
rect 283286 52808 283342 52864
rect 283194 52536 283250 52592
rect 283838 121352 283894 121408
rect 283654 118632 283710 118688
rect 283562 117000 283618 117056
rect 283746 112648 283802 112704
rect 283838 103944 283894 104000
rect 283654 99592 283710 99648
rect 283838 97996 283840 98016
rect 283840 97996 283892 98016
rect 283892 97996 283894 98016
rect 283838 97960 283894 97996
rect 283746 96600 283802 96656
rect 283654 81912 283710 81968
rect 283654 80552 283710 80608
rect 283838 95260 283894 95296
rect 283838 95240 283840 95260
rect 283840 95240 283892 95260
rect 283892 95240 283894 95260
rect 283838 93608 283894 93664
rect 283838 89256 283894 89312
rect 283838 87896 283894 87952
rect 283838 86264 283894 86320
rect 283838 68856 283894 68912
rect 283838 64504 283894 64560
rect 283838 61512 283894 61568
rect 283838 58520 283894 58576
rect 283838 46824 283894 46880
rect 283838 45464 283894 45520
rect 284206 182824 284262 182880
rect 284206 177112 284262 177168
rect 284206 174120 284262 174176
rect 284206 171148 284262 171184
rect 284206 171128 284208 171148
rect 284208 171128 284260 171148
rect 284260 171128 284262 171148
rect 284022 153720 284078 153776
rect 284206 142060 284208 142080
rect 284208 142060 284260 142080
rect 284260 142060 284262 142080
rect 284206 142024 284262 142060
rect 284206 136040 284262 136096
rect 284022 109656 284078 109712
rect 284022 108296 284078 108352
rect 284022 106936 284078 106992
rect 284206 100952 284262 101008
rect 284022 90888 284078 90944
rect 284206 78920 284262 78976
rect 284206 74588 284262 74624
rect 284206 74568 284208 74588
rect 284208 74568 284260 74588
rect 284260 74568 284262 74588
rect 284206 71848 284262 71904
rect 285218 263880 285274 263936
rect 285034 41928 285090 41984
rect 285954 37848 286010 37904
rect 287978 266872 288034 266928
rect 294602 42744 294658 42800
rect 293222 42336 293278 42392
rect 299662 569880 299718 569936
rect 299570 560360 299626 560416
rect 299294 549208 299350 549264
rect 299478 549208 299534 549264
rect 299662 521600 299718 521656
rect 299846 521600 299902 521656
rect 299478 502288 299534 502344
rect 299754 502324 299756 502344
rect 299756 502324 299808 502344
rect 299808 502324 299810 502344
rect 299754 502288 299810 502324
rect 299478 492632 299534 492688
rect 299662 492652 299718 492688
rect 299662 492632 299664 492652
rect 299664 492632 299716 492652
rect 299716 492632 299718 492652
rect 299478 412664 299534 412720
rect 299754 412664 299810 412720
rect 299202 391992 299258 392048
rect 299386 391992 299442 392048
rect 299662 273264 299718 273320
rect 299662 270544 299718 270600
rect 299478 251232 299534 251288
rect 299754 251232 299810 251288
rect 299478 241440 299534 241496
rect 299662 241440 299718 241496
rect 299478 222128 299534 222184
rect 299662 222128 299718 222184
rect 299478 183504 299534 183560
rect 299662 183504 299718 183560
rect 299478 154536 299534 154592
rect 299754 154536 299810 154592
rect 299478 135224 299534 135280
rect 299754 135224 299810 135280
rect 299478 115912 299534 115968
rect 299754 115912 299810 115968
rect 365074 686024 365130 686080
rect 364522 685888 364578 685944
rect 364154 579672 364210 579728
rect 364338 579672 364394 579728
rect 322202 267144 322258 267200
rect 364430 540912 364486 540968
rect 364614 540912 364670 540968
rect 364430 521600 364486 521656
rect 364614 521600 364670 521656
rect 364246 502288 364302 502344
rect 364522 502324 364524 502344
rect 364524 502324 364576 502344
rect 364576 502324 364578 502344
rect 364522 502288 364578 502324
rect 364246 492632 364302 492688
rect 364430 492632 364486 492688
rect 364522 268368 364578 268424
rect 356702 266464 356758 266520
rect 330022 3168 330078 3224
rect 340694 3984 340750 4040
rect 378138 29688 378194 29744
rect 393318 21256 393374 21312
rect 424874 556416 424930 556472
rect 425058 556416 425114 556472
rect 415398 556316 415400 556336
rect 415400 556316 415452 556336
rect 415452 556316 415454 556336
rect 415398 556280 415454 556316
rect 425058 555872 425114 555928
rect 429382 521600 429438 521656
rect 429566 521600 429622 521656
rect 429198 502288 429254 502344
rect 429474 502324 429476 502344
rect 429476 502324 429528 502344
rect 429528 502324 429530 502344
rect 429474 502288 429530 502324
rect 429198 492632 429254 492688
rect 429382 492652 429438 492688
rect 429382 492632 429384 492652
rect 429384 492632 429436 492652
rect 429436 492632 429438 492652
rect 429198 454008 429254 454064
rect 429474 454008 429530 454064
rect 429014 434696 429070 434752
rect 429198 434696 429254 434752
rect 429014 415384 429070 415440
rect 429198 415384 429254 415440
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 493874 579672 493930 579728
rect 494058 579672 494114 579728
rect 521658 556436 521714 556472
rect 521658 556416 521660 556436
rect 521660 556416 521712 556436
rect 521712 556416 521714 556436
rect 494150 540912 494206 540968
rect 494334 540912 494390 540968
rect 494150 521600 494206 521656
rect 494334 521600 494390 521656
rect 493966 502288 494022 502344
rect 494242 502324 494244 502344
rect 494244 502324 494296 502344
rect 494296 502324 494298 502344
rect 494242 502288 494298 502324
rect 493966 492632 494022 492688
rect 494150 492632 494206 492688
rect 529294 556144 529350 556200
rect 407762 267824 407818 267880
rect 399482 42472 399538 42528
rect 397826 9016 397882 9072
rect 401322 6840 401378 6896
rect 415398 33768 415454 33824
rect 429106 86944 429162 87000
rect 429290 86944 429346 87000
rect 429290 67496 429346 67552
rect 429566 67496 429622 67552
rect 429198 35128 429254 35184
rect 450174 3712 450230 3768
rect 454866 8880 454922 8936
rect 457258 3576 457314 3632
rect 473358 25608 473414 25664
rect 471978 25472 472034 25528
rect 487158 269184 487214 269240
rect 480258 29552 480314 29608
rect 486974 3440 487030 3496
rect 494058 266600 494114 266656
rect 511998 265376 512054 265432
rect 504822 3304 504878 3360
rect 512090 36488 512146 36544
rect 528558 265240 528614 265296
rect 526258 6704 526314 6760
rect 525062 4800 525118 4856
rect 531318 264152 531374 264208
rect 529938 32544 529994 32600
rect 580170 697992 580226 698048
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 580170 580760 580226 580816
rect 534078 556552 534134 556608
rect 540978 556552 541034 556608
rect 533986 556144 534042 556200
rect 553398 556416 553454 556472
rect 553306 556280 553362 556336
rect 540978 556144 541034 556200
rect 580170 545536 580226 545592
rect 580170 533840 580226 533896
rect 542542 521600 542598 521656
rect 542726 521600 542782 521656
rect 580170 510312 580226 510368
rect 542358 502288 542414 502344
rect 542634 502324 542636 502344
rect 542636 502324 542688 502344
rect 542688 502324 542690 502344
rect 542634 502288 542690 502324
rect 580170 498616 580226 498672
rect 542358 492632 542414 492688
rect 542542 492652 542598 492688
rect 542542 492632 542544 492652
rect 542544 492632 542596 492652
rect 542596 492632 542598 492652
rect 580170 486784 580226 486840
rect 580170 463392 580226 463448
rect 542358 454008 542414 454064
rect 542634 454008 542690 454064
rect 580170 451696 580226 451752
rect 580170 439864 580226 439920
rect 542174 434696 542230 434752
rect 542358 434696 542414 434752
rect 580170 416472 580226 416528
rect 542174 415384 542230 415440
rect 542358 415384 542414 415440
rect 580170 404776 580226 404832
rect 580170 392944 580226 393000
rect 580170 369552 580226 369608
rect 580170 357856 580226 357912
rect 580170 346024 580226 346080
rect 580170 322632 580226 322688
rect 579802 310800 579858 310856
rect 580170 299104 580226 299160
rect 580170 275712 580226 275768
rect 536930 3440 536986 3496
rect 542358 231784 542414 231840
rect 542358 106256 542414 106312
rect 554778 265784 554834 265840
rect 543738 264424 543794 264480
rect 542542 231820 542544 231840
rect 542544 231820 542596 231840
rect 542596 231820 542598 231840
rect 542542 231784 542598 231820
rect 542542 212472 542598 212528
rect 542726 212472 542782 212528
rect 542542 193160 542598 193216
rect 542726 193160 542782 193216
rect 542542 115932 542598 115968
rect 542542 115912 542544 115932
rect 542544 115912 542596 115932
rect 542596 115912 542598 115932
rect 542726 115912 542782 115968
rect 542634 106256 542690 106312
rect 542634 80008 542690 80064
rect 542634 77288 542690 77344
rect 542634 77152 542690 77208
rect 542542 67632 542598 67688
rect 542634 42064 542690 42120
rect 549258 15816 549314 15872
rect 565818 265512 565874 265568
rect 558366 6568 558422 6624
rect 563150 24112 563206 24168
rect 565542 6432 565598 6488
rect 574742 265104 574798 265160
rect 571338 32408 571394 32464
rect 569038 6296 569094 6352
rect 572626 6160 572682 6216
rect 581090 264288 581146 264344
rect 579802 263880 579858 263936
rect 575478 263744 575534 263800
rect 579802 252184 579858 252240
rect 580262 228792 580318 228848
rect 579894 205264 579950 205320
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579894 158344 579950 158400
rect 580170 134816 580226 134872
rect 579894 123120 579950 123176
rect 579894 87896 579950 87952
rect 579618 76200 579674 76256
rect 580170 64504 580226 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
<< metal3 >>
rect 57830 700436 57836 700500
rect 57900 700498 57906 700500
rect 170305 700498 170371 700501
rect 57900 700496 170371 700498
rect 57900 700440 170310 700496
rect 170366 700440 170371 700496
rect 57900 700438 170371 700440
rect 57900 700436 57906 700438
rect 170305 700435 170371 700438
rect 56358 700300 56364 700364
rect 56428 700362 56434 700364
rect 218973 700362 219039 700365
rect 56428 700360 219039 700362
rect 56428 700304 218978 700360
rect 219034 700304 219039 700360
rect 56428 700302 219039 700304
rect 56428 700300 56434 700302
rect 218973 700299 219039 700302
rect 267641 700362 267707 700365
rect 285622 700362 285628 700364
rect 267641 700360 285628 700362
rect 267641 700304 267646 700360
rect 267702 700304 285628 700360
rect 267641 700302 285628 700304
rect 267641 700299 267707 700302
rect 285622 700300 285628 700302
rect 285692 700300 285698 700364
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 365069 686082 365135 686085
rect 494881 686082 494947 686085
rect 364382 686080 365135 686082
rect 364382 686024 365074 686080
rect 365130 686024 365135 686080
rect 364382 686022 365135 686024
rect 364382 685946 364442 686022
rect 365069 686019 365135 686022
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 364517 685946 364583 685949
rect 364382 685944 364583 685946
rect 364382 685888 364522 685944
rect 364578 685888 364583 685944
rect 364382 685886 364583 685888
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 364517 685883 364583 685886
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3325 682274 3391 682277
rect -960 682272 3391 682274
rect -960 682216 3330 682272
rect 3386 682216 3391 682272
rect -960 682214 3391 682216
rect -960 682124 480 682214
rect 3325 682211 3391 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3325 653578 3391 653581
rect -960 653576 3391 653578
rect -960 653520 3330 653576
rect 3386 653520 3391 653576
rect -960 653518 3391 653520
rect -960 653428 480 653518
rect 3325 653515 3391 653518
rect 3325 652898 3391 652901
rect 57094 652898 57100 652900
rect 3325 652896 57100 652898
rect 3325 652840 3330 652896
rect 3386 652840 57100 652896
rect 3325 652838 57100 652840
rect 3325 652835 3391 652838
rect 57094 652836 57100 652838
rect 57164 652836 57170 652900
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 4061 624882 4127 624885
rect -960 624880 4127 624882
rect -960 624824 4066 624880
rect 4122 624824 4127 624880
rect -960 624822 4127 624824
rect -960 624732 480 624822
rect 4061 624819 4127 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 364149 579730 364215 579733
rect 364333 579730 364399 579733
rect 364149 579728 364399 579730
rect 364149 579672 364154 579728
rect 364210 579672 364338 579728
rect 364394 579672 364399 579728
rect 364149 579670 364399 579672
rect 364149 579667 364215 579670
rect 364333 579667 364399 579670
rect 493869 579730 493935 579733
rect 494053 579730 494119 579733
rect 493869 579728 494119 579730
rect 493869 579672 493874 579728
rect 493930 579672 494058 579728
rect 494114 579672 494119 579728
rect 493869 579670 494119 579672
rect 493869 579667 493935 579670
rect 494053 579667 494119 579670
rect 299657 569940 299723 569941
rect 299606 569938 299612 569940
rect 299566 569878 299612 569938
rect 299676 569936 299723 569940
rect 299718 569880 299723 569936
rect 299606 569876 299612 569878
rect 299676 569876 299723 569880
rect 299657 569875 299723 569876
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 4061 567354 4127 567357
rect -960 567352 4127 567354
rect -960 567296 4066 567352
rect 4122 567296 4127 567352
rect -960 567294 4127 567296
rect -960 567204 480 567294
rect 4061 567291 4127 567294
rect 299565 560420 299631 560421
rect 299565 560418 299612 560420
rect 299520 560416 299612 560418
rect 299520 560360 299570 560416
rect 299520 560358 299612 560360
rect 299565 560356 299612 560358
rect 299676 560356 299682 560420
rect 299565 560355 299631 560356
rect 583520 557290 584960 557380
rect 583342 557230 584960 557290
rect 534073 556610 534139 556613
rect 540973 556610 541039 556613
rect 534073 556608 541039 556610
rect 534073 556552 534078 556608
rect 534134 556552 540978 556608
rect 541034 556552 541039 556608
rect 534073 556550 541039 556552
rect 534073 556547 534139 556550
rect 540973 556547 541039 556550
rect 287102 556414 292682 556474
rect 286174 556140 286180 556204
rect 286244 556202 286250 556204
rect 287102 556202 287162 556414
rect 286244 556142 287162 556202
rect 292622 556202 292682 556414
rect 299422 556412 299428 556476
rect 299492 556474 299498 556476
rect 424869 556474 424935 556477
rect 425053 556474 425119 556477
rect 299492 556414 316050 556474
rect 299492 556412 299498 556414
rect 315990 556338 316050 556414
rect 325742 556414 335370 556474
rect 315990 556278 325618 556338
rect 299422 556202 299428 556204
rect 292622 556142 299428 556202
rect 286244 556140 286250 556142
rect 299422 556140 299428 556142
rect 299492 556140 299498 556204
rect 325558 556202 325618 556278
rect 325742 556202 325802 556414
rect 335310 556338 335370 556414
rect 345062 556414 354690 556474
rect 335310 556278 344938 556338
rect 325558 556142 325802 556202
rect 344878 556202 344938 556278
rect 345062 556202 345122 556414
rect 354630 556338 354690 556414
rect 364382 556414 374010 556474
rect 354630 556278 364258 556338
rect 344878 556142 345122 556202
rect 364198 556202 364258 556278
rect 364382 556202 364442 556414
rect 373950 556338 374010 556414
rect 383702 556414 393330 556474
rect 373950 556278 383578 556338
rect 364198 556142 364442 556202
rect 383518 556202 383578 556278
rect 383702 556202 383762 556414
rect 393270 556338 393330 556414
rect 403022 556414 412650 556474
rect 393270 556278 402898 556338
rect 383518 556142 383762 556202
rect 402838 556202 402898 556278
rect 403022 556202 403082 556414
rect 412590 556338 412650 556414
rect 424869 556472 425119 556474
rect 424869 556416 424874 556472
rect 424930 556416 425058 556472
rect 425114 556416 425119 556472
rect 424869 556414 425119 556416
rect 424869 556411 424935 556414
rect 425053 556411 425119 556414
rect 434662 556412 434668 556476
rect 434732 556474 434738 556476
rect 521653 556474 521719 556477
rect 434732 556414 451290 556474
rect 434732 556412 434738 556414
rect 415393 556338 415459 556341
rect 412590 556336 415459 556338
rect 412590 556280 415398 556336
rect 415454 556280 415459 556336
rect 412590 556278 415459 556280
rect 451230 556338 451290 556414
rect 460982 556414 470610 556474
rect 451230 556278 460858 556338
rect 415393 556275 415459 556278
rect 402838 556142 403082 556202
rect 460798 556202 460858 556278
rect 460982 556202 461042 556414
rect 470550 556338 470610 556414
rect 480302 556414 489930 556474
rect 470550 556278 480178 556338
rect 460798 556142 461042 556202
rect 480118 556202 480178 556278
rect 480302 556202 480362 556414
rect 489870 556338 489930 556414
rect 499622 556414 509250 556474
rect 489870 556278 499498 556338
rect 480118 556142 480362 556202
rect 499438 556202 499498 556278
rect 499622 556202 499682 556414
rect 509190 556338 509250 556414
rect 518942 556472 521719 556474
rect 518942 556416 521658 556472
rect 521714 556416 521719 556472
rect 518942 556414 521719 556416
rect 509190 556278 518818 556338
rect 499438 556142 499682 556202
rect 518758 556202 518818 556278
rect 518942 556202 519002 556414
rect 521653 556411 521719 556414
rect 553393 556474 553459 556477
rect 553393 556472 567210 556474
rect 553393 556416 553398 556472
rect 553454 556416 567210 556472
rect 553393 556414 567210 556416
rect 553393 556411 553459 556414
rect 553301 556338 553367 556341
rect 550590 556336 553367 556338
rect 550590 556280 553306 556336
rect 553362 556280 553367 556336
rect 550590 556278 553367 556280
rect 567150 556338 567210 556414
rect 583342 556338 583402 557230
rect 583520 557140 584960 557230
rect 567150 556278 576778 556338
rect 518758 556142 519002 556202
rect 529289 556202 529355 556205
rect 533981 556202 534047 556205
rect 529289 556200 534047 556202
rect 529289 556144 529294 556200
rect 529350 556144 533986 556200
rect 534042 556144 534047 556200
rect 529289 556142 534047 556144
rect 529289 556139 529355 556142
rect 533981 556139 534047 556142
rect 540973 556202 541039 556205
rect 550590 556202 550650 556278
rect 553301 556275 553367 556278
rect 540973 556200 550650 556202
rect 540973 556144 540978 556200
rect 541034 556144 550650 556200
rect 540973 556142 550650 556144
rect 576718 556202 576778 556278
rect 576902 556278 583402 556338
rect 576902 556202 576962 556278
rect 576718 556142 576962 556202
rect 540973 556139 541039 556142
rect 425053 555930 425119 555933
rect 434662 555930 434668 555932
rect 425053 555928 434668 555930
rect 425053 555872 425058 555928
rect 425114 555872 434668 555928
rect 425053 555870 434668 555872
rect 425053 555867 425119 555870
rect 434662 555868 434668 555870
rect 434732 555868 434738 555932
rect -960 553074 480 553164
rect 4061 553074 4127 553077
rect -960 553072 4127 553074
rect -960 553016 4066 553072
rect 4122 553016 4127 553072
rect -960 553014 4127 553016
rect -960 552924 480 553014
rect 4061 553011 4127 553014
rect 299289 549266 299355 549269
rect 299473 549266 299539 549269
rect 299289 549264 299539 549266
rect 299289 549208 299294 549264
rect 299350 549208 299478 549264
rect 299534 549208 299539 549264
rect 299289 549206 299539 549208
rect 299289 549203 299355 549206
rect 299473 549203 299539 549206
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 364425 540970 364491 540973
rect 364609 540970 364675 540973
rect 364425 540968 364675 540970
rect 364425 540912 364430 540968
rect 364486 540912 364614 540968
rect 364670 540912 364675 540968
rect 364425 540910 364675 540912
rect 364425 540907 364491 540910
rect 364609 540907 364675 540910
rect 494145 540970 494211 540973
rect 494329 540970 494395 540973
rect 494145 540968 494395 540970
rect 494145 540912 494150 540968
rect 494206 540912 494334 540968
rect 494390 540912 494395 540968
rect 494145 540910 494395 540912
rect 494145 540907 494211 540910
rect 494329 540907 494395 540910
rect -960 538658 480 538748
rect 3969 538658 4035 538661
rect -960 538656 4035 538658
rect -960 538600 3974 538656
rect 4030 538600 4035 538656
rect -960 538598 4035 538600
rect -960 538508 480 538598
rect 3969 538595 4035 538598
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 8109 531314 8175 531317
rect 8385 531314 8451 531317
rect 8109 531312 8451 531314
rect 8109 531256 8114 531312
rect 8170 531256 8390 531312
rect 8446 531256 8451 531312
rect 8109 531254 8451 531256
rect 8109 531251 8175 531254
rect 8385 531251 8451 531254
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 299657 521658 299723 521661
rect 299841 521658 299907 521661
rect 299657 521656 299907 521658
rect 299657 521600 299662 521656
rect 299718 521600 299846 521656
rect 299902 521600 299907 521656
rect 299657 521598 299907 521600
rect 299657 521595 299723 521598
rect 299841 521595 299907 521598
rect 364425 521658 364491 521661
rect 364609 521658 364675 521661
rect 364425 521656 364675 521658
rect 364425 521600 364430 521656
rect 364486 521600 364614 521656
rect 364670 521600 364675 521656
rect 364425 521598 364675 521600
rect 364425 521595 364491 521598
rect 364609 521595 364675 521598
rect 429377 521658 429443 521661
rect 429561 521658 429627 521661
rect 429377 521656 429627 521658
rect 429377 521600 429382 521656
rect 429438 521600 429566 521656
rect 429622 521600 429627 521656
rect 429377 521598 429627 521600
rect 429377 521595 429443 521598
rect 429561 521595 429627 521598
rect 494145 521658 494211 521661
rect 494329 521658 494395 521661
rect 494145 521656 494395 521658
rect 494145 521600 494150 521656
rect 494206 521600 494334 521656
rect 494390 521600 494395 521656
rect 494145 521598 494395 521600
rect 494145 521595 494211 521598
rect 494329 521595 494395 521598
rect 542537 521658 542603 521661
rect 542721 521658 542787 521661
rect 542537 521656 542787 521658
rect 542537 521600 542542 521656
rect 542598 521600 542726 521656
rect 542782 521600 542787 521656
rect 542537 521598 542787 521600
rect 542537 521595 542603 521598
rect 542721 521595 542787 521598
rect 8109 512002 8175 512005
rect 8385 512002 8451 512005
rect 8109 512000 8451 512002
rect 8109 511944 8114 512000
rect 8170 511944 8390 512000
rect 8446 511944 8451 512000
rect 8109 511942 8451 511944
rect 8109 511939 8175 511942
rect 8385 511939 8451 511942
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3877 509962 3943 509965
rect -960 509960 3943 509962
rect -960 509904 3882 509960
rect 3938 509904 3943 509960
rect -960 509902 3943 509904
rect -960 509812 480 509902
rect 3877 509899 3943 509902
rect 299473 502346 299539 502349
rect 299749 502346 299815 502349
rect 299473 502344 299815 502346
rect 299473 502288 299478 502344
rect 299534 502288 299754 502344
rect 299810 502288 299815 502344
rect 299473 502286 299815 502288
rect 299473 502283 299539 502286
rect 299749 502283 299815 502286
rect 364241 502346 364307 502349
rect 364517 502346 364583 502349
rect 364241 502344 364583 502346
rect 364241 502288 364246 502344
rect 364302 502288 364522 502344
rect 364578 502288 364583 502344
rect 364241 502286 364583 502288
rect 364241 502283 364307 502286
rect 364517 502283 364583 502286
rect 429193 502346 429259 502349
rect 429469 502346 429535 502349
rect 429193 502344 429535 502346
rect 429193 502288 429198 502344
rect 429254 502288 429474 502344
rect 429530 502288 429535 502344
rect 429193 502286 429535 502288
rect 429193 502283 429259 502286
rect 429469 502283 429535 502286
rect 493961 502346 494027 502349
rect 494237 502346 494303 502349
rect 493961 502344 494303 502346
rect 493961 502288 493966 502344
rect 494022 502288 494242 502344
rect 494298 502288 494303 502344
rect 493961 502286 494303 502288
rect 493961 502283 494027 502286
rect 494237 502283 494303 502286
rect 542353 502346 542419 502349
rect 542629 502346 542695 502349
rect 542353 502344 542695 502346
rect 542353 502288 542358 502344
rect 542414 502288 542634 502344
rect 542690 502288 542695 502344
rect 542353 502286 542695 502288
rect 542353 502283 542419 502286
rect 542629 502283 542695 502286
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 4061 495546 4127 495549
rect -960 495544 4127 495546
rect -960 495488 4066 495544
rect 4122 495488 4127 495544
rect -960 495486 4127 495488
rect -960 495396 480 495486
rect 4061 495483 4127 495486
rect 299473 492690 299539 492693
rect 299657 492690 299723 492693
rect 299473 492688 299723 492690
rect 299473 492632 299478 492688
rect 299534 492632 299662 492688
rect 299718 492632 299723 492688
rect 299473 492630 299723 492632
rect 299473 492627 299539 492630
rect 299657 492627 299723 492630
rect 364241 492690 364307 492693
rect 364425 492690 364491 492693
rect 364241 492688 364491 492690
rect 364241 492632 364246 492688
rect 364302 492632 364430 492688
rect 364486 492632 364491 492688
rect 364241 492630 364491 492632
rect 364241 492627 364307 492630
rect 364425 492627 364491 492630
rect 429193 492690 429259 492693
rect 429377 492690 429443 492693
rect 429193 492688 429443 492690
rect 429193 492632 429198 492688
rect 429254 492632 429382 492688
rect 429438 492632 429443 492688
rect 429193 492630 429443 492632
rect 429193 492627 429259 492630
rect 429377 492627 429443 492630
rect 493961 492690 494027 492693
rect 494145 492690 494211 492693
rect 493961 492688 494211 492690
rect 493961 492632 493966 492688
rect 494022 492632 494150 492688
rect 494206 492632 494211 492688
rect 493961 492630 494211 492632
rect 493961 492627 494027 492630
rect 494145 492627 494211 492630
rect 542353 492690 542419 492693
rect 542537 492690 542603 492693
rect 542353 492688 542603 492690
rect 542353 492632 542358 492688
rect 542414 492632 542542 492688
rect 542598 492632 542603 492688
rect 542353 492630 542603 492632
rect 542353 492627 542419 492630
rect 542537 492627 542603 492630
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 7925 483034 7991 483037
rect 8201 483034 8267 483037
rect 7925 483032 8267 483034
rect 7925 482976 7930 483032
rect 7986 482976 8206 483032
rect 8262 482976 8267 483032
rect 7925 482974 8267 482976
rect 7925 482971 7991 482974
rect 8201 482971 8267 482974
rect -960 481130 480 481220
rect 3325 481130 3391 481133
rect -960 481128 3391 481130
rect -960 481072 3330 481128
rect 3386 481072 3391 481128
rect -960 481070 3391 481072
rect -960 480980 480 481070
rect 3325 481067 3391 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 429193 454066 429259 454069
rect 429469 454066 429535 454069
rect 429193 454064 429535 454066
rect 429193 454008 429198 454064
rect 429254 454008 429474 454064
rect 429530 454008 429535 454064
rect 429193 454006 429535 454008
rect 429193 454003 429259 454006
rect 429469 454003 429535 454006
rect 542353 454066 542419 454069
rect 542629 454066 542695 454069
rect 542353 454064 542695 454066
rect 542353 454008 542358 454064
rect 542414 454008 542634 454064
rect 542690 454008 542695 454064
rect 542353 454006 542695 454008
rect 542353 454003 542419 454006
rect 542629 454003 542695 454006
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3785 438018 3851 438021
rect -960 438016 3851 438018
rect -960 437960 3790 438016
rect 3846 437960 3851 438016
rect -960 437958 3851 437960
rect -960 437868 480 437958
rect 3785 437955 3851 437958
rect 7833 434754 7899 434757
rect 8017 434754 8083 434757
rect 7833 434752 8083 434754
rect 7833 434696 7838 434752
rect 7894 434696 8022 434752
rect 8078 434696 8083 434752
rect 7833 434694 8083 434696
rect 7833 434691 7899 434694
rect 8017 434691 8083 434694
rect 429009 434754 429075 434757
rect 429193 434754 429259 434757
rect 429009 434752 429259 434754
rect 429009 434696 429014 434752
rect 429070 434696 429198 434752
rect 429254 434696 429259 434752
rect 429009 434694 429259 434696
rect 429009 434691 429075 434694
rect 429193 434691 429259 434694
rect 542169 434754 542235 434757
rect 542353 434754 542419 434757
rect 542169 434752 542419 434754
rect 542169 434696 542174 434752
rect 542230 434696 542358 434752
rect 542414 434696 542419 434752
rect 542169 434694 542419 434696
rect 542169 434691 542235 434694
rect 542353 434691 542419 434694
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 4061 423738 4127 423741
rect -960 423736 4127 423738
rect -960 423680 4066 423736
rect 4122 423680 4127 423736
rect -960 423678 4127 423680
rect -960 423588 480 423678
rect 4061 423675 4127 423678
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect 429009 415442 429075 415445
rect 429193 415442 429259 415445
rect 429009 415440 429259 415442
rect 429009 415384 429014 415440
rect 429070 415384 429198 415440
rect 429254 415384 429259 415440
rect 429009 415382 429259 415384
rect 429009 415379 429075 415382
rect 429193 415379 429259 415382
rect 542169 415442 542235 415445
rect 542353 415442 542419 415445
rect 542169 415440 542419 415442
rect 542169 415384 542174 415440
rect 542230 415384 542358 415440
rect 542414 415384 542419 415440
rect 542169 415382 542419 415384
rect 542169 415379 542235 415382
rect 542353 415379 542419 415382
rect 299473 412722 299539 412725
rect 299749 412722 299815 412725
rect 299473 412720 299815 412722
rect 299473 412664 299478 412720
rect 299534 412664 299754 412720
rect 299810 412664 299815 412720
rect 299473 412662 299815 412664
rect 299473 412659 299539 412662
rect 299749 412659 299815 412662
rect -960 409172 480 409412
rect 580165 404834 580231 404837
rect 583520 404834 584960 404924
rect 580165 404832 584960 404834
rect 580165 404776 580170 404832
rect 580226 404776 584960 404832
rect 580165 404774 584960 404776
rect 580165 404771 580231 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 4061 395042 4127 395045
rect -960 395040 4127 395042
rect -960 394984 4066 395040
rect 4122 394984 4127 395040
rect -960 394982 4127 394984
rect -960 394892 480 394982
rect 4061 394979 4127 394982
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 299197 392050 299263 392053
rect 299381 392050 299447 392053
rect 299197 392048 299447 392050
rect 299197 391992 299202 392048
rect 299258 391992 299386 392048
rect 299442 391992 299447 392048
rect 299197 391990 299447 391992
rect 299197 391987 299263 391990
rect 299381 391987 299447 391990
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3969 380626 4035 380629
rect -960 380624 4035 380626
rect -960 380568 3974 380624
rect 4030 380568 4035 380624
rect -960 380566 4035 380568
rect -960 380476 480 380566
rect 3969 380563 4035 380566
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 4061 366210 4127 366213
rect -960 366208 4127 366210
rect -960 366152 4066 366208
rect 4122 366152 4127 366208
rect -960 366150 4127 366152
rect -960 366060 480 366150
rect 4061 366147 4127 366150
rect 580165 357914 580231 357917
rect 583520 357914 584960 358004
rect 580165 357912 584960 357914
rect 580165 357856 580170 357912
rect 580226 357856 584960 357912
rect 580165 357854 584960 357856
rect 580165 357851 580231 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect -960 337514 480 337604
rect 4061 337514 4127 337517
rect -960 337512 4127 337514
rect -960 337456 4066 337512
rect 4122 337456 4127 337512
rect -960 337454 4127 337456
rect -960 337364 480 337454
rect 4061 337451 4127 337454
rect 583520 334236 584960 334476
rect -960 323098 480 323188
rect 3601 323098 3667 323101
rect -960 323096 3667 323098
rect -960 323040 3606 323096
rect 3662 323040 3667 323096
rect -960 323038 3667 323040
rect -960 322948 480 323038
rect 3601 323035 3667 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 579797 310858 579863 310861
rect 583520 310858 584960 310948
rect 579797 310856 584960 310858
rect 579797 310800 579802 310856
rect 579858 310800 584960 310856
rect 579797 310798 584960 310800
rect 579797 310795 579863 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 4061 308818 4127 308821
rect -960 308816 4127 308818
rect -960 308760 4066 308816
rect 4122 308760 4127 308816
rect -960 308758 4127 308760
rect -960 308668 480 308758
rect 4061 308755 4127 308758
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3141 294402 3207 294405
rect -960 294400 3207 294402
rect -960 294344 3146 294400
rect 3202 294344 3207 294400
rect -960 294342 3207 294344
rect -960 294252 480 294342
rect 3141 294339 3207 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3693 280122 3759 280125
rect -960 280120 3759 280122
rect -960 280064 3698 280120
rect 3754 280064 3759 280120
rect -960 280062 3759 280064
rect -960 279972 480 280062
rect 3693 280059 3759 280062
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 299657 273324 299723 273325
rect 299606 273322 299612 273324
rect 299566 273262 299612 273322
rect 299676 273320 299723 273324
rect 299718 273264 299723 273320
rect 299606 273260 299612 273262
rect 299676 273260 299723 273264
rect 299657 273259 299723 273260
rect 299657 270604 299723 270605
rect 299606 270540 299612 270604
rect 299676 270602 299723 270604
rect 299676 270600 299768 270602
rect 299718 270544 299768 270600
rect 299676 270542 299768 270544
rect 299676 270540 299723 270542
rect 299657 270539 299723 270540
rect 246021 269650 246087 269653
rect 280470 269650 280476 269652
rect 246021 269648 280476 269650
rect 246021 269592 246026 269648
rect 246082 269592 280476 269648
rect 246021 269590 280476 269592
rect 246021 269587 246087 269590
rect 280470 269588 280476 269590
rect 280540 269588 280546 269652
rect 244917 269514 244983 269517
rect 278814 269514 278820 269516
rect 244917 269512 278820 269514
rect 244917 269456 244922 269512
rect 244978 269456 278820 269512
rect 244917 269454 278820 269456
rect 244917 269451 244983 269454
rect 278814 269452 278820 269454
rect 278884 269452 278890 269516
rect 199469 269378 199535 269381
rect 282494 269378 282500 269380
rect 199469 269376 282500 269378
rect 199469 269320 199474 269376
rect 199530 269320 282500 269376
rect 199469 269318 282500 269320
rect 199469 269315 199535 269318
rect 282494 269316 282500 269318
rect 282564 269316 282570 269380
rect 74901 269242 74967 269245
rect 487153 269242 487219 269245
rect 74901 269240 487219 269242
rect 74901 269184 74906 269240
rect 74962 269184 487158 269240
rect 487214 269184 487219 269240
rect 74901 269182 487219 269184
rect 74901 269179 74967 269182
rect 487153 269179 487219 269182
rect 86677 268426 86743 268429
rect 364517 268426 364583 268429
rect 86677 268424 364583 268426
rect 86677 268368 86682 268424
rect 86738 268368 364522 268424
rect 364578 268368 364583 268424
rect 86677 268366 364583 268368
rect 86677 268363 86743 268366
rect 364517 268363 364583 268366
rect 200389 268018 200455 268021
rect 281758 268018 281764 268020
rect 200389 268016 281764 268018
rect 200389 267960 200394 268016
rect 200450 267960 281764 268016
rect 200389 267958 281764 267960
rect 200389 267955 200455 267958
rect 281758 267956 281764 267958
rect 281828 267956 281834 268020
rect 102501 267882 102567 267885
rect 407757 267882 407823 267885
rect 102501 267880 407823 267882
rect 102501 267824 102506 267880
rect 102562 267824 407762 267880
rect 407818 267824 407823 267880
rect 102501 267822 407823 267824
rect 102501 267819 102567 267822
rect 407757 267819 407823 267822
rect 280102 267548 280108 267612
rect 280172 267610 280178 267612
rect 289670 267610 289676 267612
rect 280172 267550 289676 267610
rect 280172 267548 280178 267550
rect 289670 267548 289676 267550
rect 289740 267548 289746 267612
rect 292062 267548 292068 267612
rect 292132 267610 292138 267612
rect 294638 267610 294644 267612
rect 292132 267550 294644 267610
rect 292132 267548 292138 267550
rect 294638 267548 294644 267550
rect 294708 267548 294714 267612
rect 241462 267276 241468 267340
rect 241532 267338 241538 267340
rect 244590 267338 244596 267340
rect 241532 267278 244596 267338
rect 241532 267276 241538 267278
rect 244590 267276 244596 267278
rect 244660 267276 244666 267340
rect 264789 267338 264855 267341
rect 278630 267338 278636 267340
rect 264789 267336 278636 267338
rect 264789 267280 264794 267336
rect 264850 267280 278636 267336
rect 264789 267278 278636 267280
rect 264789 267275 264855 267278
rect 278630 267276 278636 267278
rect 278700 267276 278706 267340
rect 78765 267202 78831 267205
rect 322197 267202 322263 267205
rect 78765 267200 322263 267202
rect 78765 267144 78770 267200
rect 78826 267144 322202 267200
rect 322258 267144 322263 267200
rect 78765 267142 322263 267144
rect 78765 267139 78831 267142
rect 322197 267139 322263 267142
rect 238109 267066 238175 267069
rect 281073 267066 281139 267069
rect 238109 267064 281139 267066
rect 238109 267008 238114 267064
rect 238170 267008 281078 267064
rect 281134 267008 281139 267064
rect 238109 267006 281139 267008
rect 238109 267003 238175 267006
rect 281073 267003 281139 267006
rect 107469 266932 107535 266933
rect 107469 266930 107516 266932
rect 107424 266928 107516 266930
rect 107424 266872 107474 266928
rect 107424 266870 107516 266872
rect 107469 266868 107516 266870
rect 107580 266868 107586 266932
rect 149053 266930 149119 266933
rect 287973 266930 288039 266933
rect 149053 266928 288039 266930
rect 149053 266872 149058 266928
rect 149114 266872 287978 266928
rect 288034 266872 288039 266928
rect 149053 266870 288039 266872
rect 107469 266867 107535 266868
rect 149053 266867 149119 266870
rect 287973 266867 288039 266870
rect 299422 266868 299428 266932
rect 299492 266930 299498 266932
rect 308990 266930 308996 266932
rect 299492 266870 308996 266930
rect 299492 266868 299498 266870
rect 308990 266868 308996 266870
rect 309060 266868 309066 266932
rect 320950 266868 320956 266932
rect 321020 266930 321026 266932
rect 328310 266930 328316 266932
rect 321020 266870 328316 266930
rect 321020 266868 321026 266870
rect 328310 266868 328316 266870
rect 328380 266868 328386 266932
rect 338062 266868 338068 266932
rect 338132 266930 338138 266932
rect 347630 266930 347636 266932
rect 338132 266870 347636 266930
rect 338132 266868 338138 266870
rect 347630 266868 347636 266870
rect 347700 266868 347706 266932
rect 357382 266868 357388 266932
rect 357452 266930 357458 266932
rect 366950 266930 366956 266932
rect 357452 266870 366956 266930
rect 357452 266868 357458 266870
rect 366950 266868 366956 266870
rect 367020 266868 367026 266932
rect 376886 266868 376892 266932
rect 376956 266930 376962 266932
rect 386270 266930 386276 266932
rect 376956 266870 386276 266930
rect 376956 266868 376962 266870
rect 386270 266868 386276 266870
rect 386340 266868 386346 266932
rect 396022 266868 396028 266932
rect 396092 266930 396098 266932
rect 405590 266930 405596 266932
rect 396092 266870 405596 266930
rect 396092 266868 396098 266870
rect 405590 266868 405596 266870
rect 405660 266868 405666 266932
rect 417550 266868 417556 266932
rect 417620 266930 417626 266932
rect 424910 266930 424916 266932
rect 417620 266870 424916 266930
rect 417620 266868 417626 266870
rect 424910 266868 424916 266870
rect 424980 266868 424986 266932
rect 436870 266868 436876 266932
rect 436940 266930 436946 266932
rect 444230 266930 444236 266932
rect 436940 266870 444236 266930
rect 436940 266868 436946 266870
rect 444230 266868 444236 266870
rect 444300 266868 444306 266932
rect 456190 266868 456196 266932
rect 456260 266930 456266 266932
rect 463550 266930 463556 266932
rect 456260 266870 463556 266930
rect 456260 266868 456266 266870
rect 463550 266868 463556 266870
rect 463620 266868 463626 266932
rect 475510 266868 475516 266932
rect 475580 266930 475586 266932
rect 482870 266930 482876 266932
rect 475580 266870 482876 266930
rect 475580 266868 475586 266870
rect 482870 266868 482876 266870
rect 482940 266868 482946 266932
rect 492806 266868 492812 266932
rect 492876 266930 492882 266932
rect 502190 266930 502196 266932
rect 492876 266870 502196 266930
rect 492876 266868 492882 266870
rect 502190 266868 502196 266870
rect 502260 266868 502266 266932
rect 511942 266868 511948 266932
rect 512012 266930 512018 266932
rect 521510 266930 521516 266932
rect 512012 266870 521516 266930
rect 512012 266868 512018 266870
rect 521510 266868 521516 266870
rect 521580 266868 521586 266932
rect 533838 266868 533844 266932
rect 533908 266930 533914 266932
rect 536782 266930 536788 266932
rect 533908 266870 536788 266930
rect 533908 266868 533914 266870
rect 536782 266868 536788 266870
rect 536852 266868 536858 266932
rect 103605 266794 103671 266797
rect 281257 266794 281323 266797
rect 103605 266792 281323 266794
rect 103605 266736 103610 266792
rect 103666 266736 281262 266792
rect 281318 266736 281323 266792
rect 103605 266734 281323 266736
rect 103605 266731 103671 266734
rect 281257 266731 281323 266734
rect 142061 266658 142127 266661
rect 263593 266658 263659 266661
rect 142061 266656 263659 266658
rect 142061 266600 142066 266656
rect 142122 266600 263598 266656
rect 263654 266600 263659 266656
rect 142061 266598 263659 266600
rect 142061 266595 142127 266598
rect 263593 266595 263659 266598
rect 270493 266658 270559 266661
rect 494053 266658 494119 266661
rect 270493 266656 494119 266658
rect 270493 266600 270498 266656
rect 270554 266600 494058 266656
rect 494114 266600 494119 266656
rect 270493 266598 494119 266600
rect 270493 266595 270559 266598
rect 494053 266595 494119 266598
rect 64638 266460 64644 266524
rect 64708 266522 64714 266524
rect 106549 266522 106615 266525
rect 64708 266520 106615 266522
rect 64708 266464 106554 266520
rect 106610 266464 106615 266520
rect 64708 266462 106615 266464
rect 64708 266460 64714 266462
rect 106549 266459 106615 266462
rect 129181 266522 129247 266525
rect 356697 266522 356763 266525
rect 129181 266520 356763 266522
rect 129181 266464 129186 266520
rect 129242 266464 356702 266520
rect 356758 266464 356763 266520
rect 129181 266462 356763 266464
rect 129181 266459 129247 266462
rect 356697 266459 356763 266462
rect 257797 266386 257863 266389
rect 271781 266386 271847 266389
rect 257797 266384 271847 266386
rect 257797 266328 257802 266384
rect 257858 266328 271786 266384
rect 271842 266328 271847 266384
rect 257797 266326 271847 266328
rect 257797 266323 257863 266326
rect 271781 266323 271847 266326
rect 231894 266188 231900 266252
rect 231964 266250 231970 266252
rect 241278 266250 241284 266252
rect 231964 266190 241284 266250
rect 231964 266188 231970 266190
rect 241278 266188 241284 266190
rect 241348 266188 241354 266252
rect 88701 265842 88767 265845
rect 554773 265842 554839 265845
rect 88701 265840 554839 265842
rect -960 265706 480 265796
rect 88701 265784 88706 265840
rect 88762 265784 554778 265840
rect 554834 265784 554839 265840
rect 88701 265782 554839 265784
rect 88701 265779 88767 265782
rect 554773 265779 554839 265782
rect 3877 265706 3943 265709
rect -960 265704 3943 265706
rect -960 265648 3882 265704
rect 3938 265648 3943 265704
rect -960 265646 3943 265648
rect -960 265556 480 265646
rect 3877 265643 3943 265646
rect 241053 265706 241119 265709
rect 280654 265706 280660 265708
rect 241053 265704 280660 265706
rect 241053 265648 241058 265704
rect 241114 265648 280660 265704
rect 241053 265646 280660 265648
rect 241053 265643 241119 265646
rect 280654 265644 280660 265646
rect 280724 265644 280730 265708
rect 126973 265570 127039 265573
rect 565813 265570 565879 265573
rect 126973 265568 565879 265570
rect 126973 265512 126978 265568
rect 127034 265512 565818 265568
rect 565874 265512 565879 265568
rect 126973 265510 565879 265512
rect 126973 265507 127039 265510
rect 565813 265507 565879 265510
rect 64965 265434 65031 265437
rect 511993 265434 512059 265437
rect 64965 265432 512059 265434
rect 64965 265376 64970 265432
rect 65026 265376 511998 265432
rect 512054 265376 512059 265432
rect 64965 265374 512059 265376
rect 64965 265371 65031 265374
rect 511993 265371 512059 265374
rect 79869 265298 79935 265301
rect 528553 265298 528619 265301
rect 79869 265296 528619 265298
rect 79869 265240 79874 265296
rect 79930 265240 528558 265296
rect 528614 265240 528619 265296
rect 79869 265238 528619 265240
rect 79869 265235 79935 265238
rect 528553 265235 528619 265238
rect 114461 265162 114527 265165
rect 574737 265162 574803 265165
rect 114461 265160 574803 265162
rect 114461 265104 114466 265160
rect 114522 265104 574742 265160
rect 574798 265104 574803 265160
rect 114461 265102 574803 265104
rect 114461 265099 114527 265102
rect 574737 265099 574803 265102
rect 271781 265026 271847 265029
rect 280838 265026 280844 265028
rect 271781 265024 280844 265026
rect 271781 264968 271786 265024
rect 271842 264968 280844 265024
rect 271781 264966 280844 264968
rect 271781 264963 271847 264966
rect 280838 264964 280844 264966
rect 280908 264964 280914 265028
rect 268285 264618 268351 264621
rect 279877 264618 279943 264621
rect 268285 264616 279943 264618
rect 268285 264560 268290 264616
rect 268346 264560 279882 264616
rect 279938 264560 279943 264616
rect 268285 264558 279943 264560
rect 268285 264555 268351 264558
rect 279877 264555 279943 264558
rect 209681 264482 209747 264485
rect 543733 264482 543799 264485
rect 209681 264480 543799 264482
rect 209681 264424 209686 264480
rect 209742 264424 543738 264480
rect 543794 264424 543799 264480
rect 209681 264422 543799 264424
rect 209681 264419 209747 264422
rect 543733 264419 543799 264422
rect 63217 264346 63283 264349
rect 64454 264346 64460 264348
rect 63217 264344 64460 264346
rect 63217 264288 63222 264344
rect 63278 264288 64460 264344
rect 63217 264286 64460 264288
rect 63217 264283 63283 264286
rect 64454 264284 64460 264286
rect 64524 264284 64530 264348
rect 113541 264346 113607 264349
rect 113541 264344 113650 264346
rect 113541 264288 113546 264344
rect 113602 264288 113650 264344
rect 113541 264283 113650 264288
rect 155902 264284 155908 264348
rect 155972 264346 155978 264348
rect 159541 264346 159607 264349
rect 155972 264344 159607 264346
rect 155972 264288 159546 264344
rect 159602 264288 159607 264344
rect 155972 264286 159607 264288
rect 155972 264284 155978 264286
rect 159541 264283 159607 264286
rect 163405 264346 163471 264349
rect 201677 264348 201743 264349
rect 163405 264344 163514 264346
rect 163405 264288 163410 264344
rect 163466 264288 163514 264344
rect 163405 264283 163514 264288
rect 201677 264344 201724 264348
rect 201788 264346 201794 264348
rect 222561 264346 222627 264349
rect 224902 264346 224908 264348
rect 201677 264288 201682 264344
rect 201677 264284 201724 264288
rect 201788 264286 201834 264346
rect 222561 264344 224908 264346
rect 222561 264288 222566 264344
rect 222622 264288 224908 264344
rect 222561 264286 224908 264288
rect 201788 264284 201794 264286
rect 201677 264283 201743 264284
rect 222561 264283 222627 264286
rect 224902 264284 224908 264286
rect 224972 264284 224978 264348
rect 255129 264346 255195 264349
rect 259126 264346 259132 264348
rect 255129 264344 259132 264346
rect 255129 264288 255134 264344
rect 255190 264288 259132 264344
rect 255129 264286 259132 264288
rect 255129 264283 255195 264286
rect 259126 264284 259132 264286
rect 259196 264284 259202 264348
rect 259453 264346 259519 264349
rect 268285 264346 268351 264349
rect 259453 264344 268351 264346
rect 259453 264288 259458 264344
rect 259514 264288 268290 264344
rect 268346 264288 268351 264344
rect 259453 264286 268351 264288
rect 259453 264283 259519 264286
rect 268285 264283 268351 264286
rect 275001 264346 275067 264349
rect 279366 264346 279372 264348
rect 275001 264344 279372 264346
rect 275001 264288 275006 264344
rect 275062 264288 279372 264344
rect 275001 264286 279372 264288
rect 275001 264283 275067 264286
rect 279366 264284 279372 264286
rect 279436 264284 279442 264348
rect 279877 264346 279943 264349
rect 581085 264346 581151 264349
rect 279877 264344 581151 264346
rect 279877 264288 279882 264344
rect 279938 264288 581090 264344
rect 581146 264288 581151 264344
rect 279877 264286 581151 264288
rect 279877 264283 279943 264286
rect 581085 264283 581151 264286
rect 113590 263938 113650 264283
rect 163454 264210 163514 264283
rect 531313 264210 531379 264213
rect 163454 264208 531379 264210
rect 163454 264152 531318 264208
rect 531374 264152 531379 264208
rect 163454 264150 531379 264152
rect 531313 264147 531379 264150
rect 224902 264012 224908 264076
rect 224972 264074 224978 264076
rect 281022 264074 281028 264076
rect 224972 264014 281028 264074
rect 224972 264012 224978 264014
rect 281022 264012 281028 264014
rect 281092 264012 281098 264076
rect 285213 263938 285279 263941
rect 113590 263936 285279 263938
rect 113590 263880 285218 263936
rect 285274 263880 285279 263936
rect 113590 263878 285279 263880
rect 285213 263875 285279 263878
rect 579797 263938 579863 263941
rect 583520 263938 584960 264028
rect 579797 263936 584960 263938
rect 579797 263880 579802 263936
rect 579858 263880 584960 263936
rect 579797 263878 584960 263880
rect 579797 263875 579863 263878
rect 259126 263740 259132 263804
rect 259196 263802 259202 263804
rect 575473 263802 575539 263805
rect 259196 263800 575539 263802
rect 259196 263744 575478 263800
rect 575534 263744 575539 263800
rect 583520 263788 584960 263878
rect 259196 263742 575539 263744
rect 259196 263740 259202 263742
rect 575473 263739 575539 263742
rect 63350 263604 63356 263668
rect 63420 263666 63426 263668
rect 155902 263666 155908 263668
rect 63420 263606 155908 263666
rect 63420 263604 63426 263606
rect 155902 263604 155908 263606
rect 155972 263604 155978 263668
rect 278630 263468 278636 263532
rect 278700 263530 278706 263532
rect 280981 263530 281047 263533
rect 278700 263528 281047 263530
rect 278700 263472 280986 263528
rect 281042 263472 281047 263528
rect 278700 263470 281047 263472
rect 278700 263468 278706 263470
rect 280981 263467 281047 263470
rect 283189 261762 283255 261765
rect 281612 261760 283255 261762
rect 281612 261704 283194 261760
rect 283250 261704 283255 261760
rect 281612 261702 283255 261704
rect 283189 261699 283255 261702
rect 59353 260402 59419 260405
rect 59353 260400 62100 260402
rect 59353 260344 59358 260400
rect 59414 260344 62100 260400
rect 59353 260342 62100 260344
rect 59353 260339 59419 260342
rect 60457 257410 60523 257413
rect 60457 257408 62100 257410
rect 60457 257352 60462 257408
rect 60518 257352 62100 257408
rect 60457 257350 62100 257352
rect 60457 257347 60523 257350
rect 282862 256050 282868 256052
rect 281612 255990 282868 256050
rect 282862 255988 282868 255990
rect 282932 255988 282938 256052
rect 60733 253058 60799 253061
rect 283097 253058 283163 253061
rect 60733 253056 62100 253058
rect 60733 253000 60738 253056
rect 60794 253000 62100 253056
rect 60733 252998 62100 253000
rect 281612 253056 283163 253058
rect 281612 253000 283102 253056
rect 283158 253000 283163 253056
rect 281612 252998 283163 253000
rect 60733 252995 60799 252998
rect 283097 252995 283163 252998
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect 61009 251698 61075 251701
rect 284109 251698 284175 251701
rect 61009 251696 62100 251698
rect 61009 251640 61014 251696
rect 61070 251640 62100 251696
rect 61009 251638 62100 251640
rect 281612 251696 284175 251698
rect 281612 251640 284114 251696
rect 284170 251640 284175 251696
rect 281612 251638 284175 251640
rect 61009 251635 61075 251638
rect 284109 251635 284175 251638
rect -960 251290 480 251380
rect 4061 251290 4127 251293
rect -960 251288 4127 251290
rect -960 251232 4066 251288
rect 4122 251232 4127 251288
rect -960 251230 4127 251232
rect -960 251140 480 251230
rect 4061 251227 4127 251230
rect 299473 251290 299539 251293
rect 299749 251290 299815 251293
rect 299473 251288 299815 251290
rect 299473 251232 299478 251288
rect 299534 251232 299754 251288
rect 299810 251232 299815 251288
rect 299473 251230 299815 251232
rect 299473 251227 299539 251230
rect 299749 251227 299815 251230
rect 60825 250066 60891 250069
rect 284201 250066 284267 250069
rect 60825 250064 62100 250066
rect 60825 250008 60830 250064
rect 60886 250008 62100 250064
rect 60825 250006 62100 250008
rect 281612 250064 284267 250066
rect 281612 250008 284206 250064
rect 284262 250008 284267 250064
rect 281612 250006 284267 250008
rect 60825 250003 60891 250006
rect 284201 250003 284267 250006
rect 61101 248706 61167 248709
rect 284201 248706 284267 248709
rect 61101 248704 62100 248706
rect 61101 248648 61106 248704
rect 61162 248648 62100 248704
rect 61101 248646 62100 248648
rect 281612 248704 284267 248706
rect 281612 248648 284206 248704
rect 284262 248648 284267 248704
rect 281612 248646 284267 248648
rect 61101 248643 61167 248646
rect 284201 248643 284267 248646
rect 282126 248372 282132 248436
rect 282196 248434 282202 248436
rect 283598 248434 283604 248436
rect 282196 248374 283604 248434
rect 282196 248372 282202 248374
rect 283598 248372 283604 248374
rect 283668 248372 283674 248436
rect 60774 247284 60780 247348
rect 60844 247346 60850 247348
rect 60844 247286 62100 247346
rect 60844 247284 60850 247286
rect 284201 245714 284267 245717
rect 281612 245712 284267 245714
rect 281612 245656 284206 245712
rect 284262 245656 284267 245712
rect 281612 245654 284267 245656
rect 284201 245651 284267 245654
rect 284201 244354 284267 244357
rect 281612 244352 284267 244354
rect 62622 243812 62682 244324
rect 281612 244296 284206 244352
rect 284262 244296 284267 244352
rect 281612 244294 284267 244296
rect 284201 244291 284267 244294
rect 283230 244156 283236 244220
rect 283300 244218 283306 244220
rect 283598 244218 283604 244220
rect 283300 244158 283604 244218
rect 283300 244156 283306 244158
rect 283598 244156 283604 244158
rect 283668 244156 283674 244220
rect 62614 243748 62620 243812
rect 62684 243748 62690 243812
rect 283230 241436 283236 241500
rect 283300 241498 283306 241500
rect 283557 241498 283623 241501
rect 283300 241496 283623 241498
rect 283300 241440 283562 241496
rect 283618 241440 283623 241496
rect 283300 241438 283623 241440
rect 283300 241436 283306 241438
rect 283557 241435 283623 241438
rect 299473 241498 299539 241501
rect 299657 241498 299723 241501
rect 299473 241496 299723 241498
rect 299473 241440 299478 241496
rect 299534 241440 299662 241496
rect 299718 241440 299723 241496
rect 299473 241438 299723 241440
rect 299473 241435 299539 241438
rect 299657 241435 299723 241438
rect 283189 241362 283255 241365
rect 281612 241360 283255 241362
rect 281612 241304 283194 241360
rect 283250 241304 283255 241360
rect 281612 241302 283255 241304
rect 283189 241299 283255 241302
rect 583520 240396 584960 240636
rect 59261 240002 59327 240005
rect 59261 240000 62100 240002
rect 59261 239944 59266 240000
rect 59322 239944 62100 240000
rect 59261 239942 62100 239944
rect 59261 239939 59327 239942
rect 60917 238370 60983 238373
rect 283833 238370 283899 238373
rect 60917 238368 62100 238370
rect 60917 238312 60922 238368
rect 60978 238312 62100 238368
rect 60917 238310 62100 238312
rect 281612 238368 283899 238370
rect 281612 238312 283838 238368
rect 283894 238312 283899 238368
rect 281612 238310 283899 238312
rect 60917 238307 60983 238310
rect 283833 238307 283899 238310
rect -960 237010 480 237100
rect 4061 237010 4127 237013
rect -960 237008 4127 237010
rect -960 236952 4066 237008
rect 4122 236952 4127 237008
rect -960 236950 4127 236952
rect -960 236860 480 236950
rect 4061 236947 4127 236950
rect 60457 237010 60523 237013
rect 60457 237008 62100 237010
rect 60457 236952 60462 237008
rect 60518 236952 62100 237008
rect 60457 236950 62100 236952
rect 60457 236947 60523 236950
rect 282913 235650 282979 235653
rect 281612 235648 282979 235650
rect 281612 235592 282918 235648
rect 282974 235592 282979 235648
rect 281612 235590 282979 235592
rect 282913 235587 282979 235590
rect 283833 234834 283899 234837
rect 283966 234834 283972 234836
rect 283833 234832 283972 234834
rect 283833 234776 283838 234832
rect 283894 234776 283972 234832
rect 283833 234774 283972 234776
rect 283833 234771 283899 234774
rect 283966 234772 283972 234774
rect 284036 234772 284042 234836
rect 59169 234018 59235 234021
rect 284201 234018 284267 234021
rect 59169 234016 62100 234018
rect 59169 233960 59174 234016
rect 59230 233960 62100 234016
rect 59169 233958 62100 233960
rect 281612 234016 284267 234018
rect 281612 233960 284206 234016
rect 284262 233960 284267 234016
rect 281612 233958 284267 233960
rect 59169 233955 59235 233958
rect 284201 233955 284267 233958
rect 283833 232116 283899 232117
rect 283782 232114 283788 232116
rect 283742 232054 283788 232114
rect 283852 232112 283899 232116
rect 283894 232056 283899 232112
rect 283782 232052 283788 232054
rect 283852 232052 283899 232056
rect 283833 232051 283899 232052
rect 283557 231980 283623 231981
rect 283557 231978 283604 231980
rect 283512 231976 283604 231978
rect 283512 231920 283562 231976
rect 283512 231918 283604 231920
rect 283557 231916 283604 231918
rect 283668 231916 283674 231980
rect 283557 231915 283623 231916
rect 542353 231842 542419 231845
rect 542537 231842 542603 231845
rect 542353 231840 542603 231842
rect 542353 231784 542358 231840
rect 542414 231784 542542 231840
rect 542598 231784 542603 231840
rect 542353 231782 542603 231784
rect 542353 231779 542419 231782
rect 542537 231779 542603 231782
rect 59077 229666 59143 229669
rect 59077 229664 62100 229666
rect 59077 229608 59082 229664
rect 59138 229608 62100 229664
rect 59077 229606 62100 229608
rect 59077 229603 59143 229606
rect 580257 228850 580323 228853
rect 583520 228850 584960 228940
rect 580257 228848 584960 228850
rect 580257 228792 580262 228848
rect 580318 228792 584960 228848
rect 580257 228790 584960 228792
rect 580257 228787 580323 228790
rect 583520 228700 584960 228790
rect 59670 228244 59676 228308
rect 59740 228306 59746 228308
rect 284109 228306 284175 228309
rect 59740 228246 62100 228306
rect 281612 228304 284175 228306
rect 281612 228248 284114 228304
rect 284170 228248 284175 228304
rect 281612 228246 284175 228248
rect 59740 228244 59746 228246
rect 284109 228243 284175 228246
rect 284201 226674 284267 226677
rect 281612 226672 284267 226674
rect 281612 226616 284206 226672
rect 284262 226616 284267 226672
rect 281612 226614 284267 226616
rect 284201 226611 284267 226614
rect 284201 225314 284267 225317
rect 281612 225312 284267 225314
rect 281612 225256 284206 225312
rect 284262 225256 284267 225312
rect 281612 225254 284267 225256
rect 284201 225251 284267 225254
rect 61285 223954 61351 223957
rect 61285 223952 62100 223954
rect 61285 223896 61290 223952
rect 61346 223896 62100 223952
rect 61285 223894 62100 223896
rect 61285 223891 61351 223894
rect -960 222594 480 222684
rect 2957 222594 3023 222597
rect -960 222592 3023 222594
rect -960 222536 2962 222592
rect 3018 222536 3023 222592
rect -960 222534 3023 222536
rect -960 222444 480 222534
rect 2957 222531 3023 222534
rect 59353 222322 59419 222325
rect 59353 222320 62100 222322
rect 59353 222264 59358 222320
rect 59414 222264 62100 222320
rect 59353 222262 62100 222264
rect 59353 222259 59419 222262
rect 299473 222186 299539 222189
rect 299657 222186 299723 222189
rect 299473 222184 299723 222186
rect 299473 222128 299478 222184
rect 299534 222128 299662 222184
rect 299718 222128 299723 222184
rect 299473 222126 299723 222128
rect 299473 222123 299539 222126
rect 299657 222123 299723 222126
rect 283414 221444 283420 221508
rect 283484 221444 283490 221508
rect 283422 221236 283482 221444
rect 283414 221172 283420 221236
rect 283484 221172 283490 221236
rect 59353 220962 59419 220965
rect 59353 220960 62100 220962
rect 59353 220904 59358 220960
rect 59414 220904 62100 220960
rect 59353 220902 62100 220904
rect 59353 220899 59419 220902
rect 283230 220084 283236 220148
rect 283300 220146 283306 220148
rect 283598 220146 283604 220148
rect 283300 220086 283604 220146
rect 283300 220084 283306 220086
rect 283598 220084 283604 220086
rect 283668 220084 283674 220148
rect 60917 219602 60983 219605
rect 60917 219600 62100 219602
rect 60917 219544 60922 219600
rect 60978 219544 62100 219600
rect 60917 219542 62100 219544
rect 60917 219539 60983 219542
rect 281030 219330 281090 219572
rect 281165 219330 281231 219333
rect 281030 219328 281231 219330
rect 281030 219272 281170 219328
rect 281226 219272 281231 219328
rect 281030 219270 281231 219272
rect 281165 219267 281231 219270
rect 59445 217970 59511 217973
rect 284201 217970 284267 217973
rect 59445 217968 62100 217970
rect 59445 217912 59450 217968
rect 59506 217912 62100 217968
rect 59445 217910 62100 217912
rect 281612 217968 284267 217970
rect 281612 217912 284206 217968
rect 284262 217912 284267 217968
rect 281612 217910 284267 217912
rect 59445 217907 59511 217910
rect 284201 217907 284267 217910
rect 580758 216956 580764 217020
rect 580828 217018 580834 217020
rect 583520 217018 584960 217108
rect 580828 216958 584960 217018
rect 580828 216956 580834 216958
rect 583520 216868 584960 216958
rect 59353 216610 59419 216613
rect 284201 216610 284267 216613
rect 59353 216608 62100 216610
rect 59353 216552 59358 216608
rect 59414 216552 62100 216608
rect 59353 216550 62100 216552
rect 281612 216608 284267 216610
rect 281612 216552 284206 216608
rect 284262 216552 284267 216608
rect 281612 216550 284267 216552
rect 59353 216547 59419 216550
rect 284201 216547 284267 216550
rect 59353 214978 59419 214981
rect 59353 214976 62100 214978
rect 59353 214920 59358 214976
rect 59414 214920 62100 214976
rect 59353 214918 62100 214920
rect 59353 214915 59419 214918
rect 281582 214436 281642 214948
rect 281574 214372 281580 214436
rect 281644 214372 281650 214436
rect 59353 213618 59419 213621
rect 284201 213618 284267 213621
rect 59353 213616 62100 213618
rect 59353 213560 59358 213616
rect 59414 213560 62100 213616
rect 59353 213558 62100 213560
rect 281612 213616 284267 213618
rect 281612 213560 284206 213616
rect 284262 213560 284267 213616
rect 281612 213558 284267 213560
rect 59353 213555 59419 213558
rect 284201 213555 284267 213558
rect 542537 212530 542603 212533
rect 542721 212530 542787 212533
rect 542537 212528 542787 212530
rect 542537 212472 542542 212528
rect 542598 212472 542726 212528
rect 542782 212472 542787 212528
rect 542537 212470 542787 212472
rect 542537 212467 542603 212470
rect 542721 212467 542787 212470
rect 56174 212196 56180 212260
rect 56244 212258 56250 212260
rect 284201 212258 284267 212261
rect 56244 212198 62100 212258
rect 281612 212256 284267 212258
rect 281612 212200 284206 212256
rect 284262 212200 284267 212256
rect 281612 212198 284267 212200
rect 56244 212196 56250 212198
rect 284201 212195 284267 212198
rect 60590 210564 60596 210628
rect 60660 210626 60666 210628
rect 60660 210566 62100 210626
rect 60660 210564 60666 210566
rect 283005 209676 283071 209677
rect 283005 209674 283052 209676
rect 282960 209672 283052 209674
rect 282960 209616 283010 209672
rect 282960 209614 283052 209616
rect 283005 209612 283052 209614
rect 283116 209612 283122 209676
rect 283005 209611 283071 209612
rect 283598 209402 283604 209404
rect 281582 209342 283604 209402
rect 281582 209236 281642 209342
rect 283598 209340 283604 209342
rect 283668 209340 283674 209404
rect 283414 209204 283420 209268
rect 283484 209204 283490 209268
rect 283422 208996 283482 209204
rect 283414 208932 283420 208996
rect 283484 208932 283490 208996
rect 61101 208314 61167 208317
rect 61878 208314 61884 208316
rect -960 208178 480 208268
rect 614 208254 61026 208314
rect 614 208178 674 208254
rect -960 208118 674 208178
rect -960 208028 480 208118
rect 60966 208042 61026 208254
rect 61101 208312 61884 208314
rect 61101 208256 61106 208312
rect 61162 208256 61884 208312
rect 61101 208254 61884 208256
rect 61101 208251 61167 208254
rect 61878 208252 61884 208254
rect 61948 208252 61954 208316
rect 61694 208042 61700 208044
rect 60966 207982 61700 208042
rect 61694 207980 61700 207982
rect 61764 207980 61770 208044
rect 284109 207906 284175 207909
rect 281612 207904 284175 207906
rect 281612 207848 284114 207904
rect 284170 207848 284175 207904
rect 281612 207846 284175 207848
rect 284109 207843 284175 207846
rect 59353 206274 59419 206277
rect 59353 206272 62100 206274
rect 59353 206216 59358 206272
rect 59414 206216 62100 206272
rect 59353 206214 62100 206216
rect 59353 206211 59419 206214
rect 283230 206212 283236 206276
rect 283300 206274 283306 206276
rect 283966 206274 283972 206276
rect 283300 206214 283972 206274
rect 283300 206212 283306 206214
rect 283966 206212 283972 206214
rect 284036 206212 284042 206276
rect 62389 205866 62455 205869
rect 62614 205866 62620 205868
rect 62389 205864 62620 205866
rect 62389 205808 62394 205864
rect 62450 205808 62620 205864
rect 62389 205806 62620 205808
rect 62389 205803 62455 205806
rect 62614 205804 62620 205806
rect 62684 205804 62690 205868
rect 579889 205322 579955 205325
rect 583520 205322 584960 205412
rect 579889 205320 584960 205322
rect 579889 205264 579894 205320
rect 579950 205264 584960 205320
rect 579889 205262 584960 205264
rect 579889 205259 579955 205262
rect 583520 205172 584960 205262
rect 284201 204914 284267 204917
rect 281612 204912 284267 204914
rect 281612 204856 284206 204912
rect 284262 204856 284267 204912
rect 281612 204854 284267 204856
rect 284201 204851 284267 204854
rect 59353 203282 59419 203285
rect 59353 203280 62100 203282
rect 59353 203224 59358 203280
rect 59414 203224 62100 203280
rect 59353 203222 62100 203224
rect 59353 203219 59419 203222
rect 284201 201922 284267 201925
rect 281612 201920 284267 201922
rect 281612 201864 284206 201920
rect 284262 201864 284267 201920
rect 281612 201862 284267 201864
rect 284201 201859 284267 201862
rect 62389 201514 62455 201517
rect 62614 201514 62620 201516
rect 62389 201512 62620 201514
rect 62389 201456 62394 201512
rect 62450 201456 62620 201512
rect 62389 201454 62620 201456
rect 62389 201451 62455 201454
rect 62614 201452 62620 201454
rect 62684 201452 62690 201516
rect 59118 200500 59124 200564
rect 59188 200562 59194 200564
rect 59188 200502 62100 200562
rect 59188 200500 59194 200502
rect 59353 198930 59419 198933
rect 284201 198930 284267 198933
rect 59353 198928 62100 198930
rect 59353 198872 59358 198928
rect 59414 198872 62100 198928
rect 59353 198870 62100 198872
rect 281612 198928 284267 198930
rect 281612 198872 284206 198928
rect 284262 198872 284267 198928
rect 281612 198870 284267 198872
rect 59353 198867 59419 198870
rect 284201 198867 284267 198870
rect 283557 197570 283623 197573
rect 281612 197568 283623 197570
rect 281612 197512 283562 197568
rect 283618 197512 283623 197568
rect 281612 197510 283623 197512
rect 283557 197507 283623 197510
rect 4889 194578 4955 194581
rect 12341 194578 12407 194581
rect 4889 194576 12407 194578
rect 4889 194520 4894 194576
rect 4950 194520 12346 194576
rect 12402 194520 12407 194576
rect 4889 194518 12407 194520
rect 4889 194515 4955 194518
rect 12341 194515 12407 194518
rect 22185 194578 22251 194581
rect 27613 194578 27679 194581
rect 59353 194578 59419 194581
rect 284201 194578 284267 194581
rect 22185 194576 27679 194578
rect 22185 194520 22190 194576
rect 22246 194520 27618 194576
rect 27674 194520 27679 194576
rect 22185 194518 27679 194520
rect 22185 194515 22251 194518
rect 27613 194515 27679 194518
rect 55078 194518 58082 194578
rect 12525 194442 12591 194445
rect 22001 194442 22067 194445
rect 55078 194442 55138 194518
rect 12525 194440 22067 194442
rect 12525 194384 12530 194440
rect 12586 194384 22006 194440
rect 22062 194384 22067 194440
rect 12525 194382 22067 194384
rect 12525 194379 12591 194382
rect 22001 194379 22067 194382
rect 45510 194382 55138 194442
rect 37181 194306 37247 194309
rect 45510 194306 45570 194382
rect 37181 194304 45570 194306
rect 37181 194248 37186 194304
rect 37242 194248 45570 194304
rect 37181 194246 45570 194248
rect 58022 194306 58082 194518
rect 59353 194576 62100 194578
rect 59353 194520 59358 194576
rect 59414 194520 62100 194576
rect 59353 194518 62100 194520
rect 281612 194576 284267 194578
rect 281612 194520 284206 194576
rect 284262 194520 284267 194576
rect 281612 194518 284267 194520
rect 59353 194515 59419 194518
rect 284201 194515 284267 194518
rect 60958 194306 60964 194308
rect 58022 194246 60964 194306
rect 37181 194243 37247 194246
rect 60958 194244 60964 194246
rect 61028 194244 61034 194308
rect -960 193898 480 193988
rect 4889 193898 4955 193901
rect -960 193896 4955 193898
rect -960 193840 4894 193896
rect 4950 193840 4955 193896
rect -960 193838 4955 193840
rect -960 193748 480 193838
rect 4889 193835 4955 193838
rect 583520 193476 584960 193716
rect 61285 193354 61351 193357
rect 61694 193354 61700 193356
rect 61285 193352 61700 193354
rect 61285 193296 61290 193352
rect 61346 193296 61700 193352
rect 61285 193294 61700 193296
rect 61285 193291 61351 193294
rect 61694 193292 61700 193294
rect 61764 193292 61770 193356
rect 60365 193218 60431 193221
rect 283005 193218 283071 193221
rect 60365 193216 62100 193218
rect 60365 193160 60370 193216
rect 60426 193160 62100 193216
rect 60365 193158 62100 193160
rect 281612 193216 283071 193218
rect 281612 193160 283010 193216
rect 283066 193160 283071 193216
rect 281612 193158 283071 193160
rect 60365 193155 60431 193158
rect 283005 193155 283071 193158
rect 542537 193218 542603 193221
rect 542721 193218 542787 193221
rect 542537 193216 542787 193218
rect 542537 193160 542542 193216
rect 542598 193160 542726 193216
rect 542782 193160 542787 193216
rect 542537 193158 542787 193160
rect 542537 193155 542603 193158
rect 542721 193155 542787 193158
rect 283833 192538 283899 192541
rect 283966 192538 283972 192540
rect 283833 192536 283972 192538
rect 283833 192480 283838 192536
rect 283894 192480 283972 192536
rect 283833 192478 283972 192480
rect 283833 192475 283899 192478
rect 283966 192476 283972 192478
rect 284036 192476 284042 192540
rect 61285 191586 61351 191589
rect 283465 191586 283531 191589
rect 61285 191584 62100 191586
rect 61285 191528 61290 191584
rect 61346 191528 62100 191584
rect 61285 191526 62100 191528
rect 281612 191584 283531 191586
rect 281612 191528 283470 191584
rect 283526 191528 283531 191584
rect 281612 191526 283531 191528
rect 61285 191523 61351 191526
rect 283465 191523 283531 191526
rect 60273 190226 60339 190229
rect 60273 190224 62100 190226
rect 60273 190168 60278 190224
rect 60334 190168 62100 190224
rect 60273 190166 62100 190168
rect 60273 190163 60339 190166
rect 281214 189685 281274 190196
rect 281165 189680 281274 189685
rect 281165 189624 281170 189680
rect 281226 189624 281274 189680
rect 281165 189622 281274 189624
rect 281165 189619 281231 189622
rect 59353 188866 59419 188869
rect 284201 188866 284267 188869
rect 59353 188864 62100 188866
rect 59353 188808 59358 188864
rect 59414 188808 62100 188864
rect 59353 188806 62100 188808
rect 281612 188864 284267 188866
rect 281612 188808 284206 188864
rect 284262 188808 284267 188864
rect 281612 188806 284267 188808
rect 59353 188803 59419 188806
rect 284201 188803 284267 188806
rect 58893 187234 58959 187237
rect 58893 187232 62100 187234
rect 58893 187176 58898 187232
rect 58954 187176 62100 187232
rect 58893 187174 62100 187176
rect 58893 187171 58959 187174
rect 58985 185874 59051 185877
rect 281993 185874 282059 185877
rect 58985 185872 62100 185874
rect 58985 185816 58990 185872
rect 59046 185816 62100 185872
rect 58985 185814 62100 185816
rect 281612 185872 282059 185874
rect 281612 185816 281998 185872
rect 282054 185816 282059 185872
rect 281612 185814 282059 185816
rect 58985 185811 59051 185814
rect 281993 185811 282059 185814
rect 283925 184514 283991 184517
rect 281612 184512 283991 184514
rect 281612 184456 283930 184512
rect 283986 184456 283991 184512
rect 281612 184454 283991 184456
rect 283925 184451 283991 184454
rect 62614 183834 62620 183836
rect 62438 183774 62620 183834
rect 62438 183700 62498 183774
rect 62614 183772 62620 183774
rect 62684 183772 62690 183836
rect 62430 183636 62436 183700
rect 62500 183636 62506 183700
rect 299473 183562 299539 183565
rect 299657 183562 299723 183565
rect 299473 183560 299723 183562
rect 299473 183504 299478 183560
rect 299534 183504 299662 183560
rect 299718 183504 299723 183560
rect 299473 183502 299723 183504
rect 299473 183499 299539 183502
rect 299657 183499 299723 183502
rect 59905 182882 59971 182885
rect 284201 182882 284267 182885
rect 59905 182880 62100 182882
rect 59905 182824 59910 182880
rect 59966 182824 62100 182880
rect 59905 182822 62100 182824
rect 281612 182880 284267 182882
rect 281612 182824 284206 182880
rect 284262 182824 284267 182880
rect 281612 182822 284267 182824
rect 59905 182819 59971 182822
rect 284201 182819 284267 182822
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect 59353 181522 59419 181525
rect 59353 181520 62100 181522
rect 59353 181464 59358 181520
rect 59414 181464 62100 181520
rect 59353 181462 62100 181464
rect 59353 181459 59419 181462
rect 4061 180706 4127 180709
rect 61326 180706 61332 180708
rect 4061 180704 61332 180706
rect 4061 180648 4066 180704
rect 4122 180648 61332 180704
rect 4061 180646 61332 180648
rect 4061 180643 4127 180646
rect 61326 180644 61332 180646
rect 61396 180644 61402 180708
rect 283230 180372 283236 180436
rect 283300 180434 283306 180436
rect 283833 180434 283899 180437
rect 283300 180432 283899 180434
rect 283300 180376 283838 180432
rect 283894 180376 283899 180432
rect 283300 180374 283899 180376
rect 283300 180372 283306 180374
rect 283833 180371 283899 180374
rect 283281 179890 283347 179893
rect 281612 179888 283347 179890
rect 281612 179832 283286 179888
rect 283342 179832 283347 179888
rect 281612 179830 283347 179832
rect 283281 179827 283347 179830
rect -960 179482 480 179572
rect 4061 179482 4127 179485
rect -960 179480 4127 179482
rect -960 179424 4066 179480
rect 4122 179424 4127 179480
rect -960 179422 4127 179424
rect -960 179332 480 179422
rect 4061 179419 4127 179422
rect 284201 177170 284267 177173
rect 281612 177168 284267 177170
rect 281612 177112 284206 177168
rect 284262 177112 284267 177168
rect 281612 177110 284267 177112
rect 284201 177107 284267 177110
rect 59537 175538 59603 175541
rect 59537 175536 62100 175538
rect 59537 175480 59542 175536
rect 59598 175480 62100 175536
rect 59537 175478 62100 175480
rect 59537 175475 59603 175478
rect 283230 174524 283236 174588
rect 283300 174586 283306 174588
rect 283782 174586 283788 174588
rect 283300 174526 283788 174586
rect 283300 174524 283306 174526
rect 283782 174524 283788 174526
rect 283852 174524 283858 174588
rect 58801 174178 58867 174181
rect 284201 174178 284267 174181
rect 58801 174176 62100 174178
rect 58801 174120 58806 174176
rect 58862 174120 62100 174176
rect 58801 174118 62100 174120
rect 281612 174176 284267 174178
rect 281612 174120 284206 174176
rect 284262 174120 284267 174176
rect 281612 174118 284267 174120
rect 58801 174115 58867 174118
rect 284201 174115 284267 174118
rect 60641 172818 60707 172821
rect 60641 172816 62100 172818
rect 60641 172760 60646 172816
rect 60702 172760 62100 172816
rect 60641 172758 62100 172760
rect 60641 172755 60707 172758
rect 281030 172549 281090 172788
rect 280981 172544 281090 172549
rect 280981 172488 280986 172544
rect 281042 172488 281090 172544
rect 280981 172486 281090 172488
rect 280981 172483 281047 172486
rect 58750 171124 58756 171188
rect 58820 171186 58826 171188
rect 284201 171186 284267 171189
rect 58820 171126 62100 171186
rect 281612 171184 284267 171186
rect 281612 171128 284206 171184
rect 284262 171128 284267 171184
rect 281612 171126 284267 171128
rect 58820 171124 58826 171126
rect 284201 171123 284267 171126
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 59353 168194 59419 168197
rect 283414 168194 283420 168196
rect 59353 168192 62100 168194
rect 59353 168136 59358 168192
rect 59414 168136 62100 168192
rect 59353 168134 62100 168136
rect 281612 168134 283420 168194
rect 59353 168131 59419 168134
rect 283414 168132 283420 168134
rect 283484 168132 283490 168196
rect 59353 165474 59419 165477
rect 283833 165474 283899 165477
rect 59353 165472 62100 165474
rect 59353 165416 59358 165472
rect 59414 165416 62100 165472
rect 59353 165414 62100 165416
rect 281612 165472 283899 165474
rect 281612 165416 283838 165472
rect 283894 165416 283899 165472
rect 281612 165414 283899 165416
rect 59353 165411 59419 165414
rect 283833 165411 283899 165414
rect -960 165066 480 165156
rect 3325 165066 3391 165069
rect -960 165064 3391 165066
rect -960 165008 3330 165064
rect 3386 165008 3391 165064
rect -960 165006 3391 165008
rect -960 164916 480 165006
rect 3325 165003 3391 165006
rect 61101 163842 61167 163845
rect 283833 163842 283899 163845
rect 61101 163840 62100 163842
rect 61101 163784 61106 163840
rect 61162 163784 62100 163840
rect 61101 163782 62100 163784
rect 281612 163840 283899 163842
rect 281612 163784 283838 163840
rect 283894 163784 283899 163840
rect 281612 163782 283899 163784
rect 61101 163779 61167 163782
rect 283833 163779 283899 163782
rect 283782 162482 283788 162484
rect 281612 162422 283788 162482
rect 283782 162420 283788 162422
rect 283852 162420 283858 162484
rect 58934 161060 58940 161124
rect 59004 161122 59010 161124
rect 283373 161122 283439 161125
rect 59004 161062 62100 161122
rect 281612 161120 283439 161122
rect 281612 161064 283378 161120
rect 283434 161064 283439 161120
rect 281612 161062 283439 161064
rect 59004 161060 59010 161062
rect 283373 161059 283439 161062
rect 61193 159490 61259 159493
rect 61193 159488 62100 159490
rect 61193 159432 61198 159488
rect 61254 159432 62100 159488
rect 61193 159430 62100 159432
rect 61193 159427 61259 159430
rect 579889 158402 579955 158405
rect 583520 158402 584960 158492
rect 579889 158400 584960 158402
rect 579889 158344 579894 158400
rect 579950 158344 584960 158400
rect 579889 158342 584960 158344
rect 579889 158339 579955 158342
rect 583520 158252 584960 158342
rect 62622 157180 62682 158100
rect 62614 157116 62620 157180
rect 62684 157116 62690 157180
rect 283281 156498 283347 156501
rect 281612 156496 283347 156498
rect 281612 156440 283286 156496
rect 283342 156440 283347 156496
rect 281612 156438 283347 156440
rect 283281 156435 283347 156438
rect 62062 154532 62068 154596
rect 62132 154594 62138 154596
rect 62430 154594 62436 154596
rect 62132 154534 62436 154594
rect 62132 154532 62138 154534
rect 62430 154532 62436 154534
rect 62500 154532 62506 154596
rect 280981 154594 281047 154597
rect 281349 154594 281415 154597
rect 280981 154592 281415 154594
rect 280981 154536 280986 154592
rect 281042 154536 281354 154592
rect 281410 154536 281415 154592
rect 280981 154534 281415 154536
rect 280981 154531 281047 154534
rect 281349 154531 281415 154534
rect 299473 154594 299539 154597
rect 299749 154594 299815 154597
rect 299473 154592 299815 154594
rect 299473 154536 299478 154592
rect 299534 154536 299754 154592
rect 299810 154536 299815 154592
rect 299473 154534 299815 154536
rect 299473 154531 299539 154534
rect 299749 154531 299815 154534
rect 60089 153778 60155 153781
rect 284017 153778 284083 153781
rect 60089 153776 62100 153778
rect 60089 153720 60094 153776
rect 60150 153720 62100 153776
rect 60089 153718 62100 153720
rect 281612 153776 284083 153778
rect 281612 153720 284022 153776
rect 284078 153720 284083 153776
rect 281612 153718 284083 153720
rect 60089 153715 60155 153718
rect 284017 153715 284083 153718
rect 283373 152146 283439 152149
rect 281612 152144 283439 152146
rect 281612 152088 283378 152144
rect 283434 152088 283439 152144
rect 281612 152086 283439 152088
rect 283373 152083 283439 152086
rect -960 150786 480 150876
rect 3601 150786 3667 150789
rect -960 150784 3667 150786
rect -960 150728 3606 150784
rect 3662 150728 3667 150784
rect -960 150726 3667 150728
rect -960 150636 480 150726
rect 3601 150723 3667 150726
rect 59353 150786 59419 150789
rect 59353 150784 62100 150786
rect 59353 150728 59358 150784
rect 59414 150728 62100 150784
rect 59353 150726 62100 150728
rect 59353 150723 59419 150726
rect 60549 149426 60615 149429
rect 283833 149426 283899 149429
rect 60549 149424 62100 149426
rect 60549 149368 60554 149424
rect 60610 149368 62100 149424
rect 60549 149366 62100 149368
rect 281612 149424 283899 149426
rect 281612 149368 283838 149424
rect 283894 149368 283899 149424
rect 281612 149366 283899 149368
rect 60549 149363 60615 149366
rect 283833 149363 283899 149366
rect 57646 147732 57652 147796
rect 57716 147794 57722 147796
rect 57716 147734 62100 147794
rect 57716 147732 57722 147734
rect 583520 146556 584960 146796
rect 58709 146434 58775 146437
rect 58709 146432 62100 146434
rect 58709 146376 58714 146432
rect 58770 146376 62100 146432
rect 58709 146374 62100 146376
rect 58709 146371 58775 146374
rect 58566 144740 58572 144804
rect 58636 144802 58642 144804
rect 283833 144802 283899 144805
rect 58636 144742 62100 144802
rect 281612 144800 283899 144802
rect 281612 144744 283838 144800
rect 283894 144744 283899 144800
rect 281612 144742 283899 144744
rect 58636 144740 58642 144742
rect 283833 144739 283899 144742
rect 62062 143652 62068 143716
rect 62132 143652 62138 143716
rect 62070 143578 62130 143652
rect 62614 143578 62620 143580
rect 62070 143518 62620 143578
rect 62614 143516 62620 143518
rect 62684 143516 62690 143580
rect 59353 143442 59419 143445
rect 283833 143442 283899 143445
rect 59353 143440 62100 143442
rect 59353 143384 59358 143440
rect 59414 143384 62100 143440
rect 59353 143382 62100 143384
rect 281612 143440 283899 143442
rect 281612 143384 283838 143440
rect 283894 143384 283899 143440
rect 281612 143382 283899 143384
rect 59353 143379 59419 143382
rect 283833 143379 283899 143382
rect 57329 142082 57395 142085
rect 284201 142082 284267 142085
rect 57329 142080 62100 142082
rect 57329 142024 57334 142080
rect 57390 142024 62100 142080
rect 57329 142022 62100 142024
rect 281612 142080 284267 142082
rect 281612 142024 284206 142080
rect 284262 142024 284267 142080
rect 281612 142022 284267 142024
rect 57329 142019 57395 142022
rect 284201 142019 284267 142022
rect 281214 138549 281274 139060
rect 281214 138544 281323 138549
rect 281214 138488 281262 138544
rect 281318 138488 281323 138544
rect 281214 138486 281323 138488
rect 281257 138483 281323 138486
rect 59302 137668 59308 137732
rect 59372 137730 59378 137732
rect 283741 137730 283807 137733
rect 59372 137670 62100 137730
rect 281612 137728 283807 137730
rect 281612 137672 283746 137728
rect 283802 137672 283807 137728
rect 281612 137670 283807 137672
rect 59372 137668 59378 137670
rect 283741 137667 283807 137670
rect -960 136370 480 136460
rect 3969 136370 4035 136373
rect -960 136368 4035 136370
rect -960 136312 3974 136368
rect 4030 136312 4035 136368
rect -960 136310 4035 136312
rect -960 136220 480 136310
rect 3969 136307 4035 136310
rect 284201 136098 284267 136101
rect 281612 136096 284267 136098
rect 281612 136040 284206 136096
rect 284262 136040 284267 136096
rect 281612 136038 284267 136040
rect 284201 136035 284267 136038
rect 281349 135418 281415 135421
rect 281030 135416 281415 135418
rect 281030 135360 281354 135416
rect 281410 135360 281415 135416
rect 281030 135358 281415 135360
rect 281030 135285 281090 135358
rect 281349 135355 281415 135358
rect 280981 135280 281090 135285
rect 280981 135224 280986 135280
rect 281042 135224 281090 135280
rect 280981 135222 281090 135224
rect 299473 135282 299539 135285
rect 299749 135282 299815 135285
rect 299473 135280 299815 135282
rect 299473 135224 299478 135280
rect 299534 135224 299754 135280
rect 299810 135224 299815 135280
rect 299473 135222 299815 135224
rect 280981 135219 281047 135222
rect 299473 135219 299539 135222
rect 299749 135219 299815 135222
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 60181 133106 60247 133109
rect 60181 133104 62100 133106
rect 60181 133048 60186 133104
rect 60242 133048 62100 133104
rect 60181 133046 62100 133048
rect 60181 133043 60247 133046
rect 59353 131746 59419 131749
rect 59353 131744 62100 131746
rect 59353 131688 59358 131744
rect 59414 131688 62100 131744
rect 59353 131686 62100 131688
rect 59353 131683 59419 131686
rect 59721 130386 59787 130389
rect 59721 130384 62100 130386
rect 59721 130328 59726 130384
rect 59782 130328 62100 130384
rect 59721 130326 62100 130328
rect 59721 130323 59787 130326
rect 281625 129298 281691 129301
rect 281582 129296 281691 129298
rect 281582 129240 281630 129296
rect 281686 129240 281691 129296
rect 281582 129235 281691 129240
rect 59353 128754 59419 128757
rect 59353 128752 62100 128754
rect 59353 128696 59358 128752
rect 59414 128696 62100 128752
rect 281582 128724 281642 129235
rect 59353 128694 62100 128696
rect 59353 128691 59419 128694
rect 62246 128148 62252 128212
rect 62316 128210 62322 128212
rect 62389 128210 62455 128213
rect 62316 128208 62455 128210
rect 62316 128152 62394 128208
rect 62450 128152 62455 128208
rect 62316 128150 62455 128152
rect 62316 128148 62322 128150
rect 62389 128147 62455 128150
rect 62246 128012 62252 128076
rect 62316 128074 62322 128076
rect 62614 128074 62620 128076
rect 62316 128014 62620 128074
rect 62316 128012 62322 128014
rect 62614 128012 62620 128014
rect 62684 128012 62690 128076
rect 283465 127394 283531 127397
rect 281612 127392 283531 127394
rect 281612 127336 283470 127392
rect 283526 127336 283531 127392
rect 281612 127334 283531 127336
rect 283465 127331 283531 127334
rect 282126 126924 282132 126988
rect 282196 126986 282202 126988
rect 283373 126986 283439 126989
rect 282196 126984 283439 126986
rect 282196 126928 283378 126984
rect 283434 126928 283439 126984
rect 282196 126926 283439 126928
rect 282196 126924 282202 126926
rect 283373 126923 283439 126926
rect 283373 126034 283439 126037
rect 281612 126032 283439 126034
rect 281612 125976 283378 126032
rect 283434 125976 283439 126032
rect 281612 125974 283439 125976
rect 283373 125971 283439 125974
rect 281533 124946 281599 124949
rect 281533 124944 281642 124946
rect 281533 124888 281538 124944
rect 281594 124888 281642 124944
rect 281533 124883 281642 124888
rect 281582 124372 281642 124883
rect 579889 123178 579955 123181
rect 583520 123178 584960 123268
rect 579889 123176 584960 123178
rect 579889 123120 579894 123176
rect 579950 123120 584960 123176
rect 579889 123118 584960 123120
rect 579889 123115 579955 123118
rect 60273 123042 60339 123045
rect 60273 123040 62100 123042
rect 60273 122984 60278 123040
rect 60334 122984 62100 123040
rect 583520 123028 584960 123118
rect 60273 122982 62100 122984
rect 60273 122979 60339 122982
rect -960 122090 480 122180
rect 2773 122090 2839 122093
rect -960 122088 2839 122090
rect -960 122032 2778 122088
rect 2834 122032 2839 122088
rect -960 122030 2839 122032
rect -960 121940 480 122030
rect 2773 122027 2839 122030
rect 59353 121410 59419 121413
rect 283833 121410 283899 121413
rect 59353 121408 62100 121410
rect 59353 121352 59358 121408
rect 59414 121352 62100 121408
rect 59353 121350 62100 121352
rect 281612 121408 283899 121410
rect 281612 121352 283838 121408
rect 283894 121352 283899 121408
rect 281612 121350 283899 121352
rect 59353 121347 59419 121350
rect 283833 121347 283899 121350
rect 58617 120050 58683 120053
rect 58617 120048 62100 120050
rect 58617 119992 58622 120048
rect 58678 119992 62100 120048
rect 58617 119990 62100 119992
rect 58617 119987 58683 119990
rect 59353 118690 59419 118693
rect 283649 118690 283715 118693
rect 59353 118688 62100 118690
rect 59353 118632 59358 118688
rect 59414 118632 62100 118688
rect 59353 118630 62100 118632
rect 281612 118688 283715 118690
rect 281612 118632 283654 118688
rect 283710 118632 283715 118688
rect 281612 118630 283715 118632
rect 59353 118627 59419 118630
rect 283649 118627 283715 118630
rect 62246 117268 62252 117332
rect 62316 117330 62322 117332
rect 62614 117330 62620 117332
rect 62316 117270 62620 117330
rect 62316 117268 62322 117270
rect 62614 117268 62620 117270
rect 62684 117268 62690 117332
rect 283557 117058 283623 117061
rect 281612 117056 283623 117058
rect 281612 117000 283562 117056
rect 283618 117000 283623 117056
rect 281612 116998 283623 117000
rect 283557 116995 283623 116998
rect 62389 116106 62455 116109
rect 62389 116104 62498 116106
rect 62389 116048 62394 116104
rect 62450 116048 62498 116104
rect 62389 116043 62498 116048
rect 62438 115972 62498 116043
rect 62430 115908 62436 115972
rect 62500 115908 62506 115972
rect 299473 115970 299539 115973
rect 299749 115970 299815 115973
rect 299473 115968 299815 115970
rect 299473 115912 299478 115968
rect 299534 115912 299754 115968
rect 299810 115912 299815 115968
rect 299473 115910 299815 115912
rect 299473 115907 299539 115910
rect 299749 115907 299815 115910
rect 542537 115970 542603 115973
rect 542721 115970 542787 115973
rect 542537 115968 542787 115970
rect 542537 115912 542542 115968
rect 542598 115912 542726 115968
rect 542782 115912 542787 115968
rect 542537 115910 542787 115912
rect 542537 115907 542603 115910
rect 542721 115907 542787 115910
rect 59629 112706 59695 112709
rect 283741 112706 283807 112709
rect 59629 112704 62100 112706
rect 59629 112648 59634 112704
rect 59690 112648 62100 112704
rect 59629 112646 62100 112648
rect 281612 112704 283807 112706
rect 281612 112648 283746 112704
rect 283802 112648 283807 112704
rect 281612 112646 283807 112648
rect 59629 112643 59695 112646
rect 283741 112643 283807 112646
rect 62389 111482 62455 111485
rect 62614 111482 62620 111484
rect 62389 111480 62620 111482
rect 62389 111424 62394 111480
rect 62450 111424 62620 111480
rect 62389 111422 62620 111424
rect 62389 111419 62455 111422
rect 62614 111420 62620 111422
rect 62684 111420 62690 111484
rect 580390 111420 580396 111484
rect 580460 111482 580466 111484
rect 583520 111482 584960 111572
rect 580460 111422 584960 111482
rect 580460 111420 580466 111422
rect 60641 111346 60707 111349
rect 60641 111344 62100 111346
rect 60641 111288 60646 111344
rect 60702 111288 62100 111344
rect 583520 111332 584960 111422
rect 60641 111286 62100 111288
rect 60641 111283 60707 111286
rect 60038 109652 60044 109716
rect 60108 109714 60114 109716
rect 284017 109714 284083 109717
rect 60108 109654 62100 109714
rect 281612 109712 284083 109714
rect 281612 109656 284022 109712
rect 284078 109656 284083 109712
rect 281612 109654 284083 109656
rect 60108 109652 60114 109654
rect 284017 109651 284083 109654
rect 284017 108354 284083 108357
rect 281612 108352 284083 108354
rect 281612 108296 284022 108352
rect 284078 108296 284083 108352
rect 281612 108294 284083 108296
rect 284017 108291 284083 108294
rect -960 107674 480 107764
rect 4061 107674 4127 107677
rect -960 107672 4127 107674
rect -960 107616 4066 107672
rect 4122 107616 4127 107672
rect -960 107614 4127 107616
rect -960 107524 480 107614
rect 4061 107611 4127 107614
rect 60641 106994 60707 106997
rect 284017 106994 284083 106997
rect 60641 106992 62100 106994
rect 60641 106936 60646 106992
rect 60702 106936 62100 106992
rect 60641 106934 62100 106936
rect 281612 106992 284083 106994
rect 281612 106936 284022 106992
rect 284078 106936 284083 106992
rect 281612 106934 284083 106936
rect 60641 106931 60707 106934
rect 284017 106931 284083 106934
rect 62389 106314 62455 106317
rect 62614 106314 62620 106316
rect 62389 106312 62620 106314
rect 62389 106256 62394 106312
rect 62450 106256 62620 106312
rect 62389 106254 62620 106256
rect 62389 106251 62455 106254
rect 62614 106252 62620 106254
rect 62684 106252 62690 106316
rect 542353 106314 542419 106317
rect 542629 106314 542695 106317
rect 542353 106312 542695 106314
rect 542353 106256 542358 106312
rect 542414 106256 542634 106312
rect 542690 106256 542695 106312
rect 542353 106254 542695 106256
rect 542353 106251 542419 106254
rect 542629 106251 542695 106254
rect 62205 106042 62271 106045
rect 62614 106042 62620 106044
rect 62205 106040 62620 106042
rect 62205 105984 62210 106040
rect 62266 105984 62620 106040
rect 62205 105982 62620 105984
rect 62205 105979 62271 105982
rect 62614 105980 62620 105982
rect 62684 105980 62690 106044
rect 60273 105362 60339 105365
rect 60273 105360 62100 105362
rect 60273 105304 60278 105360
rect 60334 105304 62100 105360
rect 60273 105302 62100 105304
rect 60273 105299 60339 105302
rect 281582 104957 281642 105332
rect 281582 104952 281691 104957
rect 281582 104896 281630 104952
rect 281686 104896 281691 104952
rect 281582 104894 281691 104896
rect 281625 104891 281691 104894
rect 59353 104002 59419 104005
rect 283833 104002 283899 104005
rect 59353 104000 62100 104002
rect 59353 103944 59358 104000
rect 59414 103944 62100 104000
rect 59353 103942 62100 103944
rect 281612 104000 283899 104002
rect 281612 103944 283838 104000
rect 283894 103944 283899 104000
rect 281612 103942 283899 103944
rect 59353 103939 59419 103942
rect 283833 103939 283899 103942
rect 59353 101010 59419 101013
rect 284201 101010 284267 101013
rect 59353 101008 62100 101010
rect 59353 100952 59358 101008
rect 59414 100952 62100 101008
rect 59353 100950 62100 100952
rect 281612 101008 284267 101010
rect 281612 100952 284206 101008
rect 284262 100952 284267 101008
rect 281612 100950 284267 100952
rect 59353 100947 59419 100950
rect 284201 100947 284267 100950
rect 283649 99650 283715 99653
rect 281612 99648 283715 99650
rect 281612 99592 283654 99648
rect 283710 99592 283715 99648
rect 583520 99636 584960 99876
rect 281612 99590 283715 99592
rect 283649 99587 283715 99590
rect 62205 98290 62271 98293
rect 62614 98290 62620 98292
rect 62205 98288 62620 98290
rect 62205 98232 62210 98288
rect 62266 98232 62620 98288
rect 62205 98230 62620 98232
rect 62205 98227 62271 98230
rect 62614 98228 62620 98230
rect 62684 98228 62690 98292
rect 61377 98018 61443 98021
rect 283833 98018 283899 98021
rect 60598 98016 61443 98018
rect 60598 97960 61382 98016
rect 61438 97960 61443 98016
rect 281612 98016 283899 98018
rect 60598 97958 61443 97960
rect 60598 97749 60658 97958
rect 61377 97955 61443 97958
rect 60549 97744 60658 97749
rect 60549 97688 60554 97744
rect 60610 97688 60658 97744
rect 60549 97686 60658 97688
rect 61377 97746 61443 97749
rect 62254 97746 62314 97988
rect 281612 97960 283838 98016
rect 283894 97960 283899 98016
rect 281612 97958 283899 97960
rect 283833 97955 283899 97958
rect 61377 97744 62314 97746
rect 61377 97688 61382 97744
rect 61438 97688 62314 97744
rect 61377 97686 62314 97688
rect 60549 97683 60615 97686
rect 61377 97683 61443 97686
rect 283741 96658 283807 96661
rect 281612 96656 283807 96658
rect 281612 96600 283746 96656
rect 283802 96600 283807 96656
rect 281612 96598 283807 96600
rect 283741 96595 283807 96598
rect 283833 95298 283899 95301
rect 281612 95296 283899 95298
rect 61193 94754 61259 94757
rect 62070 94754 62130 95268
rect 281612 95240 283838 95296
rect 283894 95240 283899 95296
rect 281612 95238 283899 95240
rect 283833 95235 283899 95238
rect 61193 94752 62130 94754
rect 61193 94696 61198 94752
rect 61254 94696 62130 94752
rect 61193 94694 62130 94696
rect 61193 94691 61259 94694
rect 62389 93802 62455 93805
rect 62614 93802 62620 93804
rect 62389 93800 62620 93802
rect 62389 93744 62394 93800
rect 62450 93744 62620 93800
rect 62389 93742 62620 93744
rect 62389 93739 62455 93742
rect 62614 93740 62620 93742
rect 62684 93740 62690 93804
rect 283833 93666 283899 93669
rect 281612 93664 283899 93666
rect 281612 93608 283838 93664
rect 283894 93608 283899 93664
rect 281612 93606 283899 93608
rect 283833 93603 283899 93606
rect -960 93258 480 93348
rect 3366 93258 3372 93260
rect -960 93198 3372 93258
rect -960 93108 480 93198
rect 3366 93196 3372 93198
rect 3436 93196 3442 93260
rect 282361 92306 282427 92309
rect 281612 92304 282427 92306
rect 281612 92248 282366 92304
rect 282422 92248 282427 92304
rect 281612 92246 282427 92248
rect 282361 92243 282427 92246
rect 59353 90946 59419 90949
rect 284017 90946 284083 90949
rect 59353 90944 62100 90946
rect 59353 90888 59358 90944
rect 59414 90888 62100 90944
rect 59353 90886 62100 90888
rect 281612 90944 284083 90946
rect 281612 90888 284022 90944
rect 284078 90888 284083 90944
rect 281612 90886 284083 90888
rect 59353 90883 59419 90886
rect 284017 90883 284083 90886
rect 283833 89314 283899 89317
rect 281612 89312 283899 89314
rect 281612 89256 283838 89312
rect 283894 89256 283899 89312
rect 281612 89254 283899 89256
rect 283833 89251 283899 89254
rect 62389 88634 62455 88637
rect 62614 88634 62620 88636
rect 62389 88632 62620 88634
rect 62389 88576 62394 88632
rect 62450 88576 62620 88632
rect 62389 88574 62620 88576
rect 62389 88571 62455 88574
rect 62614 88572 62620 88574
rect 62684 88572 62690 88636
rect 59721 87954 59787 87957
rect 283833 87954 283899 87957
rect 59721 87952 62100 87954
rect 59721 87896 59726 87952
rect 59782 87896 62100 87952
rect 59721 87894 62100 87896
rect 281612 87952 283899 87954
rect 281612 87896 283838 87952
rect 283894 87896 283899 87952
rect 281612 87894 283899 87896
rect 59721 87891 59787 87894
rect 283833 87891 283899 87894
rect 579889 87954 579955 87957
rect 583520 87954 584960 88044
rect 579889 87952 584960 87954
rect 579889 87896 579894 87952
rect 579950 87896 584960 87952
rect 579889 87894 584960 87896
rect 579889 87891 579955 87894
rect 583520 87804 584960 87894
rect 429101 87002 429167 87005
rect 429285 87002 429351 87005
rect 429101 87000 429351 87002
rect 429101 86944 429106 87000
rect 429162 86944 429290 87000
rect 429346 86944 429351 87000
rect 429101 86942 429351 86944
rect 429101 86939 429167 86942
rect 429285 86939 429351 86942
rect 61377 86322 61443 86325
rect 283833 86322 283899 86325
rect 61377 86320 62100 86322
rect 61377 86264 61382 86320
rect 61438 86264 62100 86320
rect 61377 86262 62100 86264
rect 281612 86320 283899 86322
rect 281612 86264 283838 86320
rect 283894 86264 283899 86320
rect 281612 86262 283899 86264
rect 61377 86259 61443 86262
rect 283833 86259 283899 86262
rect 281214 84421 281274 84932
rect 281165 84416 281274 84421
rect 281165 84360 281170 84416
rect 281226 84360 281274 84416
rect 281165 84358 281274 84360
rect 281165 84355 281231 84358
rect 59629 83602 59695 83605
rect 281901 83602 281967 83605
rect 59629 83600 62100 83602
rect 59629 83544 59634 83600
rect 59690 83544 62100 83600
rect 59629 83542 62100 83544
rect 281612 83600 281967 83602
rect 281612 83544 281906 83600
rect 281962 83544 281967 83600
rect 281612 83542 281967 83544
rect 59629 83539 59695 83542
rect 281901 83539 281967 83542
rect 283649 81970 283715 81973
rect 281612 81968 283715 81970
rect 62438 81565 62498 81940
rect 281612 81912 283654 81968
rect 283710 81912 283715 81968
rect 281612 81910 283715 81912
rect 283649 81907 283715 81910
rect 60181 81562 60247 81565
rect 61142 81562 61148 81564
rect 60181 81560 61148 81562
rect 60181 81504 60186 81560
rect 60242 81504 61148 81560
rect 60181 81502 61148 81504
rect 60181 81499 60247 81502
rect 61142 81500 61148 81502
rect 61212 81500 61218 81564
rect 62389 81560 62498 81565
rect 62389 81504 62394 81560
rect 62450 81504 62498 81560
rect 62389 81502 62498 81504
rect 62389 81499 62455 81502
rect 59997 80610 60063 80613
rect 283649 80610 283715 80613
rect 59997 80608 62100 80610
rect 59997 80552 60002 80608
rect 60058 80552 62100 80608
rect 59997 80550 62100 80552
rect 281612 80608 283715 80610
rect 281612 80552 283654 80608
rect 283710 80552 283715 80608
rect 281612 80550 283715 80552
rect 59997 80547 60063 80550
rect 283649 80547 283715 80550
rect 542629 80068 542695 80069
rect 542629 80064 542676 80068
rect 542740 80066 542746 80068
rect 542629 80008 542634 80064
rect 542629 80004 542676 80008
rect 542740 80006 542786 80066
rect 542740 80004 542746 80006
rect 542629 80003 542695 80004
rect 62297 79930 62363 79933
rect 62614 79930 62620 79932
rect 62297 79928 62620 79930
rect 62297 79872 62302 79928
rect 62358 79872 62620 79928
rect 62297 79870 62620 79872
rect 62297 79867 62363 79870
rect 62614 79868 62620 79870
rect 62684 79868 62690 79932
rect 19558 79188 19564 79252
rect 19628 79250 19634 79252
rect 22686 79250 22692 79252
rect 19628 79190 22692 79250
rect 19628 79188 19634 79190
rect 22686 79188 22692 79190
rect 22756 79188 22762 79252
rect 28942 79188 28948 79252
rect 29012 79250 29018 79252
rect 42006 79250 42012 79252
rect 29012 79190 42012 79250
rect 29012 79188 29018 79190
rect 42006 79188 42012 79190
rect 42076 79188 42082 79252
rect 60089 79250 60155 79253
rect 60089 79248 62100 79250
rect 60089 79192 60094 79248
rect 60150 79192 62100 79248
rect 60089 79190 62100 79192
rect 60089 79187 60155 79190
rect -960 78978 480 79068
rect 3969 78978 4035 78981
rect 284201 78978 284267 78981
rect -960 78976 4035 78978
rect -960 78920 3974 78976
rect 4030 78920 4035 78976
rect -960 78918 4035 78920
rect 281612 78976 284267 78978
rect 281612 78920 284206 78976
rect 284262 78920 284267 78976
rect 281612 78918 284267 78920
rect -960 78828 480 78918
rect 3969 78915 4035 78918
rect 284201 78915 284267 78918
rect 59353 77618 59419 77621
rect 59353 77616 62100 77618
rect 59353 77560 59358 77616
rect 59414 77560 62100 77616
rect 59353 77558 62100 77560
rect 59353 77555 59419 77558
rect 542629 77348 542695 77349
rect 542629 77344 542676 77348
rect 542740 77346 542746 77348
rect 542629 77288 542634 77344
rect 542629 77284 542676 77288
rect 542740 77286 542786 77346
rect 542740 77284 542746 77286
rect 542629 77283 542695 77284
rect 494830 77148 494836 77212
rect 494900 77210 494906 77212
rect 500718 77210 500724 77212
rect 494900 77150 500724 77210
rect 494900 77148 494906 77150
rect 500718 77148 500724 77150
rect 500788 77148 500794 77212
rect 542486 77148 542492 77212
rect 542556 77210 542562 77212
rect 542629 77210 542695 77213
rect 542556 77208 542695 77210
rect 542556 77152 542634 77208
rect 542690 77152 542695 77208
rect 542556 77150 542695 77152
rect 542556 77148 542562 77150
rect 542629 77147 542695 77150
rect 62246 76468 62252 76532
rect 62316 76468 62322 76532
rect 281390 76468 281396 76532
rect 281460 76530 281466 76532
rect 297950 76530 297956 76532
rect 281460 76470 297956 76530
rect 281460 76468 281466 76470
rect 297950 76468 297956 76470
rect 298020 76468 298026 76532
rect 376702 76468 376708 76532
rect 376772 76530 376778 76532
rect 389766 76530 389772 76532
rect 376772 76470 389772 76530
rect 376772 76468 376778 76470
rect 389766 76468 389772 76470
rect 389836 76468 389842 76532
rect 62254 76228 62314 76468
rect 282085 76258 282151 76261
rect 281612 76256 282151 76258
rect 281612 76200 282090 76256
rect 282146 76200 282151 76256
rect 281612 76198 282151 76200
rect 282085 76195 282151 76198
rect 579613 76258 579679 76261
rect 583520 76258 584960 76348
rect 579613 76256 584960 76258
rect 579613 76200 579618 76256
rect 579674 76200 584960 76256
rect 579613 76198 584960 76200
rect 579613 76195 579679 76198
rect 583520 76108 584960 76198
rect 60457 75852 60523 75853
rect 60406 75850 60412 75852
rect 60366 75790 60412 75850
rect 60476 75848 60523 75852
rect 60518 75792 60523 75848
rect 60406 75788 60412 75790
rect 60476 75788 60523 75792
rect 347814 75788 347820 75852
rect 347884 75850 347890 75852
rect 357198 75850 357204 75852
rect 347884 75790 357204 75850
rect 347884 75788 347890 75790
rect 357198 75788 357204 75790
rect 357268 75788 357274 75852
rect 60457 75787 60523 75788
rect 59353 74626 59419 74629
rect 284201 74626 284267 74629
rect 59353 74624 62100 74626
rect 59353 74568 59358 74624
rect 59414 74568 62100 74624
rect 59353 74566 62100 74568
rect 281612 74624 284267 74626
rect 281612 74568 284206 74624
rect 284262 74568 284267 74624
rect 281612 74566 284267 74568
rect 59353 74563 59419 74566
rect 284201 74563 284267 74566
rect 61009 73130 61075 73133
rect 61510 73130 61516 73132
rect 61009 73128 61516 73130
rect 61009 73072 61014 73128
rect 61070 73072 61516 73128
rect 61009 73070 61516 73072
rect 61009 73067 61075 73070
rect 61510 73068 61516 73070
rect 61580 73068 61586 73132
rect 288382 73068 288388 73132
rect 288452 73130 288458 73132
rect 297950 73130 297956 73132
rect 288452 73070 297956 73130
rect 288452 73068 288458 73070
rect 297950 73068 297956 73070
rect 298020 73068 298026 73132
rect 552606 73068 552612 73132
rect 552676 73130 552682 73132
rect 553526 73130 553532 73132
rect 552676 73070 553532 73130
rect 552676 73068 552682 73070
rect 553526 73068 553532 73070
rect 553596 73068 553602 73132
rect 281390 72388 281396 72452
rect 281460 72450 281466 72452
rect 283414 72450 283420 72452
rect 281460 72390 283420 72450
rect 281460 72388 281466 72390
rect 283414 72388 283420 72390
rect 283484 72388 283490 72452
rect 378542 72388 378548 72452
rect 378612 72450 378618 72452
rect 386270 72450 386276 72452
rect 378612 72390 386276 72450
rect 378612 72388 378618 72390
rect 386270 72388 386276 72390
rect 386340 72388 386346 72452
rect 415710 72388 415716 72452
rect 415780 72450 415786 72452
rect 424910 72450 424916 72452
rect 415780 72390 424916 72450
rect 415780 72388 415786 72390
rect 424910 72388 424916 72390
rect 424980 72388 424986 72452
rect 437238 72388 437244 72452
rect 437308 72450 437314 72452
rect 444230 72450 444236 72452
rect 437308 72390 444236 72450
rect 437308 72388 437314 72390
rect 444230 72388 444236 72390
rect 444300 72388 444306 72452
rect 475326 72388 475332 72452
rect 475396 72450 475402 72452
rect 476246 72450 476252 72452
rect 475396 72390 476252 72450
rect 475396 72388 475402 72390
rect 476246 72388 476252 72390
rect 476316 72388 476322 72452
rect 284201 71906 284267 71909
rect 281612 71904 284267 71906
rect 281612 71848 284206 71904
rect 284262 71848 284267 71904
rect 281612 71846 284267 71848
rect 284201 71843 284267 71846
rect 309174 71708 309180 71772
rect 309244 71770 309250 71772
rect 318558 71770 318564 71772
rect 309244 71710 318564 71770
rect 309244 71708 309250 71710
rect 318558 71708 318564 71710
rect 318628 71708 318634 71772
rect 328494 71708 328500 71772
rect 328564 71770 328570 71772
rect 337878 71770 337884 71772
rect 328564 71710 337884 71770
rect 328564 71708 328570 71710
rect 337878 71708 337884 71710
rect 337948 71708 337954 71772
rect 347814 71708 347820 71772
rect 347884 71770 347890 71772
rect 357198 71770 357204 71772
rect 347884 71710 357204 71770
rect 347884 71708 347890 71710
rect 357198 71708 357204 71710
rect 357268 71708 357274 71772
rect 367134 71708 367140 71772
rect 367204 71770 367210 71772
rect 376518 71770 376524 71772
rect 367204 71710 376524 71770
rect 367204 71708 367210 71710
rect 376518 71708 376524 71710
rect 376588 71708 376594 71772
rect 453982 71708 453988 71772
rect 454052 71770 454058 71772
rect 463550 71770 463556 71772
rect 454052 71710 463556 71770
rect 454052 71708 454058 71710
rect 463550 71708 463556 71710
rect 463620 71708 463626 71772
rect 502374 71708 502380 71772
rect 502444 71770 502450 71772
rect 511758 71770 511764 71772
rect 502444 71710 511764 71770
rect 502444 71708 502450 71710
rect 511758 71708 511764 71710
rect 511828 71708 511834 71772
rect 62205 70546 62271 70549
rect 62614 70546 62620 70548
rect 62205 70544 62620 70546
rect 62205 70488 62210 70544
rect 62266 70488 62620 70544
rect 62205 70486 62620 70488
rect 62205 70483 62271 70486
rect 62614 70484 62620 70486
rect 62684 70484 62690 70548
rect 61009 70274 61075 70277
rect 61009 70272 62100 70274
rect 61009 70216 61014 70272
rect 61070 70216 62100 70272
rect 61009 70214 62100 70216
rect 61009 70211 61075 70214
rect 283833 68914 283899 68917
rect 281612 68912 283899 68914
rect 281612 68856 283838 68912
rect 283894 68856 283899 68912
rect 281612 68854 283899 68856
rect 283833 68851 283899 68854
rect 62297 67826 62363 67829
rect 62614 67826 62620 67828
rect 62297 67824 62620 67826
rect 62297 67768 62302 67824
rect 62358 67768 62620 67824
rect 62297 67766 62620 67768
rect 62297 67763 62363 67766
rect 62614 67764 62620 67766
rect 62684 67764 62690 67828
rect 542537 67692 542603 67693
rect 542486 67628 542492 67692
rect 542556 67690 542603 67692
rect 542556 67688 542648 67690
rect 542598 67632 542648 67688
rect 542556 67630 542648 67632
rect 542556 67628 542603 67630
rect 542537 67627 542603 67628
rect 429285 67554 429351 67557
rect 429561 67554 429627 67557
rect 429285 67552 429627 67554
rect 429285 67496 429290 67552
rect 429346 67496 429566 67552
rect 429622 67496 429627 67552
rect 429285 67494 429627 67496
rect 429285 67491 429351 67494
rect 429561 67491 429627 67494
rect 59353 65922 59419 65925
rect 59353 65920 62100 65922
rect 59353 65864 59358 65920
rect 59414 65864 62100 65920
rect 59353 65862 62100 65864
rect 59353 65859 59419 65862
rect 281582 65381 281642 65892
rect 281533 65376 281642 65381
rect 281533 65320 281538 65376
rect 281594 65320 281642 65376
rect 281533 65318 281642 65320
rect 281533 65315 281599 65318
rect -960 64562 480 64652
rect 3509 64562 3575 64565
rect -960 64560 3575 64562
rect -960 64504 3514 64560
rect 3570 64504 3575 64560
rect -960 64502 3575 64504
rect -960 64412 480 64502
rect 3509 64499 3575 64502
rect 59905 64562 59971 64565
rect 283833 64562 283899 64565
rect 59905 64560 62100 64562
rect 59905 64504 59910 64560
rect 59966 64504 62100 64560
rect 59905 64502 62100 64504
rect 281612 64560 283899 64562
rect 281612 64504 283838 64560
rect 283894 64504 283899 64560
rect 281612 64502 283899 64504
rect 59905 64499 59971 64502
rect 283833 64499 283899 64502
rect 580165 64562 580231 64565
rect 583520 64562 584960 64652
rect 580165 64560 584960 64562
rect 580165 64504 580170 64560
rect 580226 64504 584960 64560
rect 580165 64502 584960 64504
rect 580165 64499 580231 64502
rect 583520 64412 584960 64502
rect 281901 62930 281967 62933
rect 281612 62928 281967 62930
rect 281612 62872 281906 62928
rect 281962 62872 281967 62928
rect 281612 62870 281967 62872
rect 281901 62867 281967 62870
rect 60038 61508 60044 61572
rect 60108 61570 60114 61572
rect 283833 61570 283899 61573
rect 60108 61510 62100 61570
rect 281612 61568 283899 61570
rect 281612 61512 283838 61568
rect 283894 61512 283899 61568
rect 281612 61510 283899 61512
rect 60108 61508 60114 61510
rect 283833 61507 283899 61510
rect 281073 60890 281139 60893
rect 281390 60890 281396 60892
rect 281073 60888 281396 60890
rect 281073 60832 281078 60888
rect 281134 60832 281396 60888
rect 281073 60830 281396 60832
rect 281073 60827 281139 60830
rect 281390 60828 281396 60830
rect 281460 60828 281466 60892
rect 62205 60754 62271 60757
rect 62614 60754 62620 60756
rect 62205 60752 62620 60754
rect 62205 60696 62210 60752
rect 62266 60696 62620 60752
rect 62205 60694 62620 60696
rect 62205 60691 62271 60694
rect 62614 60692 62620 60694
rect 62684 60692 62690 60756
rect 59353 60210 59419 60213
rect 59353 60208 62100 60210
rect 59353 60152 59358 60208
rect 59414 60152 62100 60208
rect 59353 60150 62100 60152
rect 59353 60147 59419 60150
rect 281030 59669 281090 60180
rect 281030 59664 281139 59669
rect 281030 59608 281078 59664
rect 281134 59608 281139 59664
rect 281030 59606 281139 59608
rect 281073 59603 281139 59606
rect 61469 58578 61535 58581
rect 283833 58578 283899 58581
rect 61469 58576 62100 58578
rect 61469 58520 61474 58576
rect 61530 58520 62100 58576
rect 61469 58518 62100 58520
rect 281612 58576 283899 58578
rect 281612 58520 283838 58576
rect 283894 58520 283899 58576
rect 281612 58518 283899 58520
rect 61469 58515 61535 58518
rect 283833 58515 283899 58518
rect 62254 53957 62314 54196
rect 62254 53952 62363 53957
rect 62254 53896 62302 53952
rect 62358 53896 62363 53952
rect 62254 53894 62363 53896
rect 62297 53891 62363 53894
rect 283281 52866 283347 52869
rect 281612 52864 283347 52866
rect 281612 52808 283286 52864
rect 283342 52808 283347 52864
rect 281612 52806 283347 52808
rect 283281 52803 283347 52806
rect 583520 52716 584960 52956
rect 283189 52596 283255 52597
rect 283189 52594 283236 52596
rect 283144 52592 283236 52594
rect 283144 52536 283194 52592
rect 283144 52534 283236 52536
rect 283189 52532 283236 52534
rect 283300 52532 283306 52596
rect 283189 52531 283255 52532
rect 62062 52396 62068 52460
rect 62132 52458 62138 52460
rect 62614 52458 62620 52460
rect 62132 52398 62620 52458
rect 62132 52396 62138 52398
rect 62614 52396 62620 52398
rect 62684 52396 62690 52460
rect 281942 52396 281948 52460
rect 282012 52458 282018 52460
rect 282821 52458 282887 52461
rect 282012 52456 282887 52458
rect 282012 52400 282826 52456
rect 282882 52400 282887 52456
rect 282012 52398 282887 52400
rect 282012 52396 282018 52398
rect 282821 52395 282887 52398
rect 282269 51234 282335 51237
rect 281612 51232 282335 51234
rect 281612 51176 282274 51232
rect 282330 51176 282335 51232
rect 281612 51174 282335 51176
rect 282269 51171 282335 51174
rect -960 50146 480 50236
rect 3509 50146 3575 50149
rect -960 50144 3575 50146
rect -960 50088 3514 50144
rect 3570 50088 3575 50144
rect -960 50086 3575 50088
rect -960 49996 480 50086
rect 3509 50083 3575 50086
rect 62070 49738 62130 49844
rect 60598 49678 62130 49738
rect 60457 49602 60523 49605
rect 60598 49602 60658 49678
rect 60457 49600 60658 49602
rect 60457 49544 60462 49600
rect 60518 49544 60658 49600
rect 60457 49542 60658 49544
rect 60457 49539 60523 49542
rect 62254 48244 62314 48484
rect 62246 48180 62252 48244
rect 62316 48180 62322 48244
rect 283833 46882 283899 46885
rect 281612 46880 283899 46882
rect 62070 46341 62130 46852
rect 281612 46824 283838 46880
rect 283894 46824 283899 46880
rect 281612 46822 283899 46824
rect 283833 46819 283899 46822
rect 62021 46336 62130 46341
rect 62021 46280 62026 46336
rect 62082 46280 62130 46336
rect 62021 46278 62130 46280
rect 62021 46275 62087 46278
rect 283833 45522 283899 45525
rect 281612 45520 283899 45522
rect 62254 44981 62314 45492
rect 281612 45464 283838 45520
rect 283894 45464 283899 45520
rect 281612 45462 283899 45464
rect 283833 45459 283899 45462
rect 62205 44976 62314 44981
rect 62205 44920 62210 44976
rect 62266 44920 62314 44976
rect 62205 44918 62314 44920
rect 62205 44915 62271 44918
rect 62246 43828 62252 43892
rect 62316 43890 62322 43892
rect 62982 43890 62988 43892
rect 62316 43830 62988 43890
rect 62316 43828 62322 43830
rect 62982 43828 62988 43830
rect 63052 43828 63058 43892
rect 63534 43828 63540 43892
rect 63604 43890 63610 43892
rect 65374 43890 65380 43892
rect 63604 43830 65380 43890
rect 63604 43828 63610 43830
rect 65374 43828 65380 43830
rect 65444 43828 65450 43892
rect 277025 43890 277091 43893
rect 277158 43890 277164 43892
rect 277025 43888 277164 43890
rect 277025 43832 277030 43888
rect 277086 43832 277164 43888
rect 277025 43830 277164 43832
rect 277025 43827 277091 43830
rect 277158 43828 277164 43830
rect 277228 43828 277234 43892
rect 62062 43692 62068 43756
rect 62132 43754 62138 43756
rect 62798 43754 62804 43756
rect 62132 43694 62804 43754
rect 62132 43692 62138 43694
rect 62798 43692 62804 43694
rect 62868 43692 62874 43756
rect 142061 43482 142127 43485
rect 281758 43482 281764 43484
rect 142061 43480 281764 43482
rect 142061 43424 142066 43480
rect 142122 43424 281764 43480
rect 142061 43422 281764 43424
rect 142061 43419 142127 43422
rect 281758 43420 281764 43422
rect 281828 43420 281834 43484
rect 79317 42802 79383 42805
rect 294597 42802 294663 42805
rect 79317 42800 294663 42802
rect 79317 42744 79322 42800
rect 79378 42744 294602 42800
rect 294658 42744 294663 42800
rect 79317 42742 294663 42744
rect 79317 42739 79383 42742
rect 294597 42739 294663 42742
rect 86309 42666 86375 42669
rect 286174 42666 286180 42668
rect 86309 42664 286180 42666
rect 86309 42608 86314 42664
rect 86370 42608 286180 42664
rect 86309 42606 286180 42608
rect 86309 42603 86375 42606
rect 286174 42604 286180 42606
rect 286244 42604 286250 42668
rect 57094 42468 57100 42532
rect 57164 42530 57170 42532
rect 158437 42530 158503 42533
rect 57164 42528 158503 42530
rect 57164 42472 158442 42528
rect 158498 42472 158503 42528
rect 57164 42470 158503 42472
rect 57164 42468 57170 42470
rect 158437 42467 158503 42470
rect 205909 42530 205975 42533
rect 399477 42530 399543 42533
rect 205909 42528 399543 42530
rect 205909 42472 205914 42528
rect 205970 42472 399482 42528
rect 399538 42472 399543 42528
rect 205909 42470 399543 42472
rect 205909 42467 205975 42470
rect 399477 42467 399543 42470
rect 161381 42394 161447 42397
rect 293217 42394 293283 42397
rect 161381 42392 293283 42394
rect 161381 42336 161386 42392
rect 161442 42336 293222 42392
rect 293278 42336 293283 42392
rect 161381 42334 293283 42336
rect 161381 42331 161447 42334
rect 293217 42331 293283 42334
rect 153101 42258 153167 42261
rect 276974 42258 276980 42260
rect 153101 42256 276980 42258
rect 153101 42200 153106 42256
rect 153162 42200 276980 42256
rect 153101 42198 276980 42200
rect 153101 42195 153167 42198
rect 276974 42196 276980 42198
rect 277044 42196 277050 42260
rect 121453 42122 121519 42125
rect 542629 42122 542695 42125
rect 121453 42120 542695 42122
rect 121453 42064 121458 42120
rect 121514 42064 542634 42120
rect 542690 42064 542695 42120
rect 121453 42062 542695 42064
rect 121453 42059 121519 42062
rect 542629 42059 542695 42062
rect 190085 41986 190151 41989
rect 285029 41986 285095 41989
rect 190085 41984 285095 41986
rect 190085 41928 190090 41984
rect 190146 41928 285034 41984
rect 285090 41928 285095 41984
rect 190085 41926 285095 41928
rect 190085 41923 190151 41926
rect 285029 41923 285095 41926
rect 56358 41244 56364 41308
rect 56428 41306 56434 41308
rect 100109 41306 100175 41309
rect 56428 41304 100175 41306
rect 56428 41248 100114 41304
rect 100170 41248 100175 41304
rect 56428 41246 100175 41248
rect 56428 41244 56434 41246
rect 100109 41243 100175 41246
rect 57830 41108 57836 41172
rect 57900 41170 57906 41172
rect 101029 41170 101095 41173
rect 57900 41168 101095 41170
rect 57900 41112 101034 41168
rect 101090 41112 101095 41168
rect 57900 41110 101095 41112
rect 57900 41108 57906 41110
rect 101029 41107 101095 41110
rect 168373 41170 168439 41173
rect 285622 41170 285628 41172
rect 168373 41168 285628 41170
rect 168373 41112 168378 41168
rect 168434 41112 285628 41168
rect 168373 41110 285628 41112
rect 168373 41107 168439 41110
rect 285622 41108 285628 41110
rect 285692 41108 285698 41172
rect 221733 41034 221799 41037
rect 283046 41034 283052 41036
rect 221733 41032 283052 41034
rect 221733 40976 221738 41032
rect 221794 40976 283052 41032
rect 221733 40974 283052 40976
rect 221733 40971 221799 40974
rect 283046 40972 283052 40974
rect 283116 40972 283122 41036
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 96061 40898 96127 40901
rect 281942 40898 281948 40900
rect 96061 40896 281948 40898
rect 96061 40840 96066 40896
rect 96122 40840 281948 40896
rect 96061 40838 281948 40840
rect 96061 40835 96127 40838
rect 281942 40836 281948 40838
rect 282012 40836 282018 40900
rect 583520 40884 584960 40974
rect 194501 39402 194567 39405
rect 278814 39402 278820 39404
rect 194501 39400 278820 39402
rect 194501 39344 194506 39400
rect 194562 39344 278820 39400
rect 194501 39342 278820 39344
rect 194501 39339 194567 39342
rect 278814 39340 278820 39342
rect 278884 39340 278890 39404
rect 136541 39266 136607 39269
rect 280470 39266 280476 39268
rect 136541 39264 280476 39266
rect 136541 39208 136546 39264
rect 136602 39208 280476 39264
rect 136541 39206 280476 39208
rect 136541 39203 136607 39206
rect 280470 39204 280476 39206
rect 280540 39204 280546 39268
rect 62430 37844 62436 37908
rect 62500 37906 62506 37908
rect 285949 37906 286015 37909
rect 62500 37904 286015 37906
rect 62500 37848 285954 37904
rect 286010 37848 286015 37904
rect 62500 37846 286015 37848
rect 62500 37844 62506 37846
rect 285949 37843 286015 37846
rect 61510 36484 61516 36548
rect 61580 36546 61586 36548
rect 512085 36546 512151 36549
rect 61580 36544 512151 36546
rect 61580 36488 512090 36544
rect 512146 36488 512151 36544
rect 61580 36486 512151 36488
rect 61580 36484 61586 36486
rect 512085 36483 512151 36486
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 61694 35124 61700 35188
rect 61764 35186 61770 35188
rect 429193 35186 429259 35189
rect 61764 35184 429259 35186
rect 61764 35128 429198 35184
rect 429254 35128 429259 35184
rect 61764 35126 429259 35128
rect 61764 35124 61770 35126
rect 429193 35123 429259 35126
rect 60590 33764 60596 33828
rect 60660 33826 60666 33828
rect 415393 33826 415459 33829
rect 60660 33824 415459 33826
rect 60660 33768 415398 33824
rect 415454 33768 415459 33824
rect 60660 33766 415459 33768
rect 60660 33764 60666 33766
rect 415393 33763 415459 33766
rect 60406 32540 60412 32604
rect 60476 32602 60482 32604
rect 529933 32602 529999 32605
rect 60476 32600 529999 32602
rect 60476 32544 529938 32600
rect 529994 32544 529999 32600
rect 60476 32542 529999 32544
rect 60476 32540 60482 32542
rect 529933 32539 529999 32542
rect 59118 32404 59124 32468
rect 59188 32466 59194 32468
rect 571333 32466 571399 32469
rect 59188 32464 571399 32466
rect 59188 32408 571338 32464
rect 571394 32408 571399 32464
rect 59188 32406 571399 32408
rect 59188 32404 59194 32406
rect 571333 32403 571399 32406
rect 64086 31860 64092 31924
rect 64156 31922 64162 31924
rect 64156 31862 64338 31922
rect 64156 31860 64162 31862
rect 64278 31788 64338 31862
rect 64270 31724 64276 31788
rect 64340 31724 64346 31788
rect 62614 30908 62620 30972
rect 62684 30970 62690 30972
rect 183553 30970 183619 30973
rect 62684 30968 183619 30970
rect 62684 30912 183558 30968
rect 183614 30912 183619 30968
rect 62684 30910 183619 30912
rect 62684 30908 62690 30910
rect 183553 30907 183619 30910
rect 139301 29882 139367 29885
rect 283230 29882 283236 29884
rect 139301 29880 283236 29882
rect 139301 29824 139306 29880
rect 139362 29824 283236 29880
rect 139301 29822 283236 29824
rect 139301 29819 139367 29822
rect 283230 29820 283236 29822
rect 283300 29820 283306 29884
rect 60774 29684 60780 29748
rect 60844 29746 60850 29748
rect 378133 29746 378199 29749
rect 60844 29744 378199 29746
rect 60844 29688 378138 29744
rect 378194 29688 378199 29744
rect 60844 29686 378199 29688
rect 60844 29684 60850 29686
rect 378133 29683 378199 29686
rect 60038 29548 60044 29612
rect 60108 29610 60114 29612
rect 480253 29610 480319 29613
rect 60108 29608 480319 29610
rect 60108 29552 480258 29608
rect 480314 29552 480319 29608
rect 60108 29550 480319 29552
rect 60108 29548 60114 29550
rect 480253 29547 480319 29550
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect 150617 29066 150683 29069
rect 150801 29066 150867 29069
rect 150617 29064 150867 29066
rect 150617 29008 150622 29064
rect 150678 29008 150806 29064
rect 150862 29008 150867 29064
rect 150617 29006 150867 29008
rect 150617 29003 150683 29006
rect 150801 29003 150867 29006
rect 64454 28188 64460 28252
rect 64524 28250 64530 28252
rect 146293 28250 146359 28253
rect 64524 28248 146359 28250
rect 64524 28192 146298 28248
rect 146354 28192 146359 28248
rect 64524 28190 146359 28192
rect 64524 28188 64530 28190
rect 146293 28187 146359 28190
rect 62982 25604 62988 25668
rect 63052 25666 63058 25668
rect 473353 25666 473419 25669
rect 63052 25664 473419 25666
rect 63052 25608 473358 25664
rect 473414 25608 473419 25664
rect 63052 25606 473419 25608
rect 63052 25604 63058 25606
rect 473353 25603 473419 25606
rect 59302 25468 59308 25532
rect 59372 25530 59378 25532
rect 471973 25530 472039 25533
rect 59372 25528 472039 25530
rect 59372 25472 471978 25528
rect 472034 25472 472039 25528
rect 59372 25470 472039 25472
rect 59372 25468 59378 25470
rect 471973 25467 472039 25470
rect 58750 24108 58756 24172
rect 58820 24170 58826 24172
rect 563145 24170 563211 24173
rect 58820 24168 563211 24170
rect 58820 24112 563150 24168
rect 563206 24112 563211 24168
rect 58820 24110 563211 24112
rect 58820 24108 58826 24110
rect 563145 24107 563211 24110
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 61878 21252 61884 21316
rect 61948 21314 61954 21316
rect 393313 21314 393379 21317
rect 61948 21312 393379 21314
rect 61948 21256 393318 21312
rect 393374 21256 393379 21312
rect 61948 21254 393379 21256
rect 61948 21252 61954 21254
rect 393313 21251 393379 21254
rect 64270 19348 64276 19412
rect 64340 19348 64346 19412
rect 64278 19140 64338 19348
rect 64270 19076 64276 19140
rect 64340 19076 64346 19140
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect 160001 16010 160067 16013
rect 282862 16010 282868 16012
rect 160001 16008 282868 16010
rect 160001 15952 160006 16008
rect 160062 15952 282868 16008
rect 160001 15950 282868 15952
rect 160001 15947 160067 15950
rect 282862 15948 282868 15950
rect 282932 15948 282938 16012
rect 58566 15812 58572 15876
rect 58636 15874 58642 15876
rect 549253 15874 549319 15877
rect 58636 15872 549319 15874
rect 58636 15816 549258 15872
rect 549314 15816 549319 15872
rect 58636 15814 549319 15816
rect 58636 15812 58642 15814
rect 549253 15811 549319 15814
rect 54753 9074 54819 9077
rect 397821 9074 397887 9077
rect 54753 9072 397887 9074
rect 54753 9016 54758 9072
rect 54814 9016 397826 9072
rect 397882 9016 397887 9072
rect 54753 9014 397887 9016
rect 54753 9011 54819 9014
rect 397821 9011 397887 9014
rect 53465 8938 53531 8941
rect 454861 8938 454927 8941
rect 53465 8936 454927 8938
rect 53465 8880 53470 8936
rect 53526 8880 454866 8936
rect 454922 8880 454927 8936
rect 53465 8878 454927 8880
rect 53465 8875 53531 8878
rect 454861 8875 454927 8878
rect -960 7170 480 7260
rect 2957 7170 3023 7173
rect -960 7168 3023 7170
rect -960 7112 2962 7168
rect 3018 7112 3023 7168
rect -960 7110 3023 7112
rect -960 7020 480 7110
rect 2957 7107 3023 7110
rect 65374 6836 65380 6900
rect 65444 6898 65450 6900
rect 172973 6898 173039 6901
rect 65444 6896 173039 6898
rect 65444 6840 172978 6896
rect 173034 6840 173039 6896
rect 65444 6838 173039 6840
rect 65444 6836 65450 6838
rect 172973 6835 173039 6838
rect 277158 6836 277164 6900
rect 277228 6898 277234 6900
rect 401317 6898 401383 6901
rect 277228 6896 401383 6898
rect 277228 6840 401322 6896
rect 401378 6840 401383 6896
rect 277228 6838 401383 6840
rect 277228 6836 277234 6838
rect 401317 6835 401383 6838
rect 55857 6762 55923 6765
rect 526253 6762 526319 6765
rect 55857 6760 526319 6762
rect 55857 6704 55862 6760
rect 55918 6704 526258 6760
rect 526314 6704 526319 6760
rect 55857 6702 526319 6704
rect 55857 6699 55923 6702
rect 526253 6699 526319 6702
rect 56174 6564 56180 6628
rect 56244 6626 56250 6628
rect 558361 6626 558427 6629
rect 56244 6624 558427 6626
rect 56244 6568 558366 6624
rect 558422 6568 558427 6624
rect 56244 6566 558427 6568
rect 56244 6564 56250 6566
rect 558361 6563 558427 6566
rect 57646 6428 57652 6492
rect 57716 6490 57722 6492
rect 565537 6490 565603 6493
rect 57716 6488 565603 6490
rect 57716 6432 565542 6488
rect 565598 6432 565603 6488
rect 57716 6430 565603 6432
rect 57716 6428 57722 6430
rect 565537 6427 565603 6430
rect 56041 6354 56107 6357
rect 569033 6354 569099 6357
rect 56041 6352 569099 6354
rect 56041 6296 56046 6352
rect 56102 6296 569038 6352
rect 569094 6296 569099 6352
rect 56041 6294 569099 6296
rect 56041 6291 56107 6294
rect 569033 6291 569099 6294
rect 57237 6218 57303 6221
rect 572621 6218 572687 6221
rect 57237 6216 572687 6218
rect 57237 6160 57242 6216
rect 57298 6160 572626 6216
rect 572682 6160 572687 6216
rect 57237 6158 572687 6160
rect 57237 6155 57303 6158
rect 572621 6155 572687 6158
rect 209865 6082 209931 6085
rect 284334 6082 284340 6084
rect 209865 6080 284340 6082
rect 209865 6024 209870 6080
rect 209926 6024 284340 6080
rect 209865 6022 284340 6024
rect 209865 6019 209931 6022
rect 284334 6020 284340 6022
rect 284404 6020 284410 6084
rect 583520 5796 584960 6036
rect 58934 4796 58940 4860
rect 59004 4858 59010 4860
rect 525057 4858 525123 4861
rect 59004 4856 525123 4858
rect 59004 4800 525062 4856
rect 525118 4800 525123 4856
rect 59004 4798 525123 4800
rect 59004 4796 59010 4798
rect 525057 4795 525123 4798
rect 56133 4042 56199 4045
rect 280061 4042 280127 4045
rect 56133 4040 280127 4042
rect 56133 3984 56138 4040
rect 56194 3984 280066 4040
rect 280122 3984 280127 4040
rect 56133 3982 280127 3984
rect 56133 3979 56199 3982
rect 280061 3979 280127 3982
rect 281022 3980 281028 4044
rect 281092 4042 281098 4044
rect 340689 4042 340755 4045
rect 281092 4040 340755 4042
rect 281092 3984 340694 4040
rect 340750 3984 340755 4040
rect 281092 3982 340755 3984
rect 281092 3980 281098 3982
rect 340689 3979 340755 3982
rect 126605 3906 126671 3909
rect 282126 3906 282132 3908
rect 126605 3904 282132 3906
rect 126605 3848 126610 3904
rect 126666 3848 282132 3904
rect 126605 3846 282132 3848
rect 126605 3843 126671 3846
rect 282126 3844 282132 3846
rect 282196 3844 282202 3908
rect 63902 3708 63908 3772
rect 63972 3770 63978 3772
rect 171777 3770 171843 3773
rect 63972 3768 171843 3770
rect 63972 3712 171782 3768
rect 171838 3712 171843 3768
rect 63972 3710 171843 3712
rect 63972 3708 63978 3710
rect 171777 3707 171843 3710
rect 280838 3708 280844 3772
rect 280908 3770 280914 3772
rect 450169 3770 450235 3773
rect 280908 3768 450235 3770
rect 280908 3712 450174 3768
rect 450230 3712 450235 3768
rect 280908 3710 450235 3712
rect 280908 3708 280914 3710
rect 450169 3707 450235 3710
rect 64638 3572 64644 3636
rect 64708 3634 64714 3636
rect 200389 3634 200455 3637
rect 64708 3632 200455 3634
rect 64708 3576 200394 3632
rect 200450 3576 200455 3632
rect 64708 3574 200455 3576
rect 64708 3572 64714 3574
rect 200389 3571 200455 3574
rect 232497 3634 232563 3637
rect 279734 3634 279740 3636
rect 232497 3632 279740 3634
rect 232497 3576 232502 3632
rect 232558 3576 279740 3632
rect 232497 3574 279740 3576
rect 232497 3571 232563 3574
rect 279734 3572 279740 3574
rect 279804 3572 279810 3636
rect 280654 3572 280660 3636
rect 280724 3634 280730 3636
rect 457253 3634 457319 3637
rect 280724 3632 457319 3634
rect 280724 3576 457258 3632
rect 457314 3576 457319 3632
rect 280724 3574 457319 3576
rect 280724 3572 280730 3574
rect 457253 3571 457319 3574
rect 57329 3498 57395 3501
rect 486969 3498 487035 3501
rect 57329 3496 487035 3498
rect 57329 3440 57334 3496
rect 57390 3440 486974 3496
rect 487030 3440 487035 3496
rect 57329 3438 487035 3440
rect 57329 3435 57395 3438
rect 486969 3435 487035 3438
rect 536782 3436 536788 3500
rect 536852 3498 536858 3500
rect 536925 3498 536991 3501
rect 536852 3496 536991 3498
rect 536852 3440 536930 3496
rect 536986 3440 536991 3496
rect 536852 3438 536991 3440
rect 536852 3436 536858 3438
rect 536925 3435 536991 3438
rect 57421 3362 57487 3365
rect 504817 3362 504883 3365
rect 57421 3360 504883 3362
rect 57421 3304 57426 3360
rect 57482 3304 504822 3360
rect 504878 3304 504883 3360
rect 57421 3302 504883 3304
rect 57421 3299 57487 3302
rect 504817 3299 504883 3302
rect 63718 3164 63724 3228
rect 63788 3226 63794 3228
rect 139669 3226 139735 3229
rect 63788 3224 139735 3226
rect 63788 3168 139674 3224
rect 139730 3168 139735 3224
rect 63788 3166 139735 3168
rect 63788 3164 63794 3166
rect 139669 3163 139735 3166
rect 279366 3164 279372 3228
rect 279436 3226 279442 3228
rect 330017 3226 330083 3229
rect 279436 3224 330083 3226
rect 279436 3168 330022 3224
rect 330078 3168 330083 3224
rect 279436 3166 330083 3168
rect 279436 3164 279442 3166
rect 330017 3163 330083 3166
<< via3 >>
rect 57836 700436 57900 700500
rect 56364 700300 56428 700364
rect 285628 700300 285692 700364
rect 57100 652836 57164 652900
rect 299612 569936 299676 569940
rect 299612 569880 299662 569936
rect 299662 569880 299676 569936
rect 299612 569876 299676 569880
rect 299612 560416 299676 560420
rect 299612 560360 299626 560416
rect 299626 560360 299676 560416
rect 299612 560356 299676 560360
rect 286180 556140 286244 556204
rect 299428 556412 299492 556476
rect 299428 556140 299492 556204
rect 434668 556412 434732 556476
rect 434668 555868 434732 555932
rect 299612 273320 299676 273324
rect 299612 273264 299662 273320
rect 299662 273264 299676 273320
rect 299612 273260 299676 273264
rect 299612 270600 299676 270604
rect 299612 270544 299662 270600
rect 299662 270544 299676 270600
rect 299612 270540 299676 270544
rect 280476 269588 280540 269652
rect 278820 269452 278884 269516
rect 282500 269316 282564 269380
rect 281764 267956 281828 268020
rect 280108 267548 280172 267612
rect 289676 267548 289740 267612
rect 292068 267548 292132 267612
rect 294644 267548 294708 267612
rect 241468 267276 241532 267340
rect 244596 267276 244660 267340
rect 278636 267276 278700 267340
rect 107516 266928 107580 266932
rect 107516 266872 107530 266928
rect 107530 266872 107580 266928
rect 107516 266868 107580 266872
rect 299428 266868 299492 266932
rect 308996 266868 309060 266932
rect 320956 266868 321020 266932
rect 328316 266868 328380 266932
rect 338068 266868 338132 266932
rect 347636 266868 347700 266932
rect 357388 266868 357452 266932
rect 366956 266868 367020 266932
rect 376892 266868 376956 266932
rect 386276 266868 386340 266932
rect 396028 266868 396092 266932
rect 405596 266868 405660 266932
rect 417556 266868 417620 266932
rect 424916 266868 424980 266932
rect 436876 266868 436940 266932
rect 444236 266868 444300 266932
rect 456196 266868 456260 266932
rect 463556 266868 463620 266932
rect 475516 266868 475580 266932
rect 482876 266868 482940 266932
rect 492812 266868 492876 266932
rect 502196 266868 502260 266932
rect 511948 266868 512012 266932
rect 521516 266868 521580 266932
rect 533844 266868 533908 266932
rect 536788 266868 536852 266932
rect 64644 266460 64708 266524
rect 231900 266188 231964 266252
rect 241284 266188 241348 266252
rect 280660 265644 280724 265708
rect 280844 264964 280908 265028
rect 64460 264284 64524 264348
rect 155908 264284 155972 264348
rect 201724 264344 201788 264348
rect 201724 264288 201738 264344
rect 201738 264288 201788 264344
rect 201724 264284 201788 264288
rect 224908 264284 224972 264348
rect 259132 264284 259196 264348
rect 279372 264284 279436 264348
rect 224908 264012 224972 264076
rect 281028 264012 281092 264076
rect 259132 263740 259196 263804
rect 63356 263604 63420 263668
rect 155908 263604 155972 263668
rect 278636 263468 278700 263532
rect 282868 255988 282932 256052
rect 282132 248372 282196 248436
rect 283604 248372 283668 248436
rect 60780 247284 60844 247348
rect 283236 244156 283300 244220
rect 283604 244156 283668 244220
rect 62620 243748 62684 243812
rect 283236 241436 283300 241500
rect 283972 234772 284036 234836
rect 283788 232112 283852 232116
rect 283788 232056 283838 232112
rect 283838 232056 283852 232112
rect 283788 232052 283852 232056
rect 283604 231976 283668 231980
rect 283604 231920 283618 231976
rect 283618 231920 283668 231976
rect 283604 231916 283668 231920
rect 59676 228244 59740 228308
rect 283420 221444 283484 221508
rect 283420 221172 283484 221236
rect 283236 220084 283300 220148
rect 283604 220084 283668 220148
rect 580764 216956 580828 217020
rect 281580 214372 281644 214436
rect 56180 212196 56244 212260
rect 60596 210564 60660 210628
rect 283052 209672 283116 209676
rect 283052 209616 283066 209672
rect 283066 209616 283116 209672
rect 283052 209612 283116 209616
rect 283604 209340 283668 209404
rect 283420 209204 283484 209268
rect 283420 208932 283484 208996
rect 61884 208252 61948 208316
rect 61700 207980 61764 208044
rect 283236 206212 283300 206276
rect 283972 206212 284036 206276
rect 62620 205804 62684 205868
rect 62620 201452 62684 201516
rect 59124 200500 59188 200564
rect 60964 194244 61028 194308
rect 61700 193292 61764 193356
rect 283972 192476 284036 192540
rect 62620 183772 62684 183836
rect 62436 183636 62500 183700
rect 61332 180644 61396 180708
rect 283236 180372 283300 180436
rect 283236 174524 283300 174588
rect 283788 174524 283852 174588
rect 58756 171124 58820 171188
rect 283420 168132 283484 168196
rect 283788 162420 283852 162484
rect 58940 161060 59004 161124
rect 62620 157116 62684 157180
rect 62068 154532 62132 154596
rect 62436 154532 62500 154596
rect 57652 147732 57716 147796
rect 58572 144740 58636 144804
rect 62068 143652 62132 143716
rect 62620 143516 62684 143580
rect 59308 137668 59372 137732
rect 62252 128148 62316 128212
rect 62252 128012 62316 128076
rect 62620 128012 62684 128076
rect 282132 126924 282196 126988
rect 62252 117268 62316 117332
rect 62620 117268 62684 117332
rect 62436 115908 62500 115972
rect 62620 111420 62684 111484
rect 580396 111420 580460 111484
rect 60044 109652 60108 109716
rect 62620 106252 62684 106316
rect 62620 105980 62684 106044
rect 62620 98228 62684 98292
rect 62620 93740 62684 93804
rect 3372 93196 3436 93260
rect 62620 88572 62684 88636
rect 61148 81500 61212 81564
rect 542676 80064 542740 80068
rect 542676 80008 542690 80064
rect 542690 80008 542740 80064
rect 542676 80004 542740 80008
rect 62620 79868 62684 79932
rect 19564 79188 19628 79252
rect 22692 79188 22756 79252
rect 28948 79188 29012 79252
rect 42012 79188 42076 79252
rect 542676 77344 542740 77348
rect 542676 77288 542690 77344
rect 542690 77288 542740 77344
rect 542676 77284 542740 77288
rect 494836 77148 494900 77212
rect 500724 77148 500788 77212
rect 542492 77148 542556 77212
rect 62252 76468 62316 76532
rect 281396 76468 281460 76532
rect 297956 76468 298020 76532
rect 376708 76468 376772 76532
rect 389772 76468 389836 76532
rect 60412 75848 60476 75852
rect 60412 75792 60462 75848
rect 60462 75792 60476 75848
rect 60412 75788 60476 75792
rect 347820 75788 347884 75852
rect 357204 75788 357268 75852
rect 61516 73068 61580 73132
rect 288388 73068 288452 73132
rect 297956 73068 298020 73132
rect 552612 73068 552676 73132
rect 553532 73068 553596 73132
rect 281396 72388 281460 72452
rect 283420 72388 283484 72452
rect 378548 72388 378612 72452
rect 386276 72388 386340 72452
rect 415716 72388 415780 72452
rect 424916 72388 424980 72452
rect 437244 72388 437308 72452
rect 444236 72388 444300 72452
rect 475332 72388 475396 72452
rect 476252 72388 476316 72452
rect 309180 71708 309244 71772
rect 318564 71708 318628 71772
rect 328500 71708 328564 71772
rect 337884 71708 337948 71772
rect 347820 71708 347884 71772
rect 357204 71708 357268 71772
rect 367140 71708 367204 71772
rect 376524 71708 376588 71772
rect 453988 71708 454052 71772
rect 463556 71708 463620 71772
rect 502380 71708 502444 71772
rect 511764 71708 511828 71772
rect 62620 70484 62684 70548
rect 62620 67764 62684 67828
rect 542492 67688 542556 67692
rect 542492 67632 542542 67688
rect 542542 67632 542556 67688
rect 542492 67628 542556 67632
rect 60044 61508 60108 61572
rect 281396 60828 281460 60892
rect 62620 60692 62684 60756
rect 283236 52592 283300 52596
rect 283236 52536 283250 52592
rect 283250 52536 283300 52592
rect 283236 52532 283300 52536
rect 62068 52396 62132 52460
rect 62620 52396 62684 52460
rect 281948 52396 282012 52460
rect 62252 48180 62316 48244
rect 62252 43828 62316 43892
rect 62988 43828 63052 43892
rect 63540 43828 63604 43892
rect 65380 43828 65444 43892
rect 277164 43828 277228 43892
rect 62068 43692 62132 43756
rect 62804 43692 62868 43756
rect 281764 43420 281828 43484
rect 286180 42604 286244 42668
rect 57100 42468 57164 42532
rect 276980 42196 277044 42260
rect 56364 41244 56428 41308
rect 57836 41108 57900 41172
rect 285628 41108 285692 41172
rect 283052 40972 283116 41036
rect 281948 40836 282012 40900
rect 278820 39340 278884 39404
rect 280476 39204 280540 39268
rect 62436 37844 62500 37908
rect 61516 36484 61580 36548
rect 61700 35124 61764 35188
rect 60596 33764 60660 33828
rect 60412 32540 60476 32604
rect 59124 32404 59188 32468
rect 64092 31860 64156 31924
rect 64276 31724 64340 31788
rect 62620 30908 62684 30972
rect 283236 29820 283300 29884
rect 60780 29684 60844 29748
rect 60044 29548 60108 29612
rect 64460 28188 64524 28252
rect 62988 25604 63052 25668
rect 59308 25468 59372 25532
rect 58756 24108 58820 24172
rect 61884 21252 61948 21316
rect 64276 19348 64340 19412
rect 64276 19076 64340 19140
rect 282868 15948 282932 16012
rect 58572 15812 58636 15876
rect 65380 6836 65444 6900
rect 277164 6836 277228 6900
rect 56180 6564 56244 6628
rect 57652 6428 57716 6492
rect 284340 6020 284404 6084
rect 58940 4796 59004 4860
rect 281028 3980 281092 4044
rect 282132 3844 282196 3908
rect 63908 3708 63972 3772
rect 280844 3708 280908 3772
rect 64644 3572 64708 3636
rect 279740 3572 279804 3636
rect 280660 3572 280724 3636
rect 536788 3436 536852 3500
rect 63724 3164 63788 3228
rect 279372 3164 279436 3228
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 -6926 -7976 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 -5986 -7036 709922
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 -5046 -6096 708982
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 -4106 -5156 708042
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 -3166 -4216 707102
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 -2226 -3276 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 3371 93260 3437 93261
rect 3371 93196 3372 93260
rect 3436 93196 3437 93260
rect 3371 93195 3437 93196
rect 3374 79338 3434 93195
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 18804 56454 19404 91898
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 19563 79252 19629 79253
rect 19563 79188 19564 79252
rect 19628 79188 19629 79252
rect 19563 79187 19629 79188
rect 19566 77978 19626 79187
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 36804 74454 37404 109898
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 57835 700500 57901 700501
rect 57835 700436 57836 700500
rect 57900 700436 57901 700500
rect 57835 700435 57901 700436
rect 56363 700364 56429 700365
rect 56363 700300 56364 700364
rect 56428 700300 56429 700364
rect 56363 700299 56429 700300
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 56179 212260 56245 212261
rect 56179 212196 56180 212260
rect 56244 212196 56245 212260
rect 56179 212195 56245 212196
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 56182 6629 56242 212195
rect 56366 41309 56426 700299
rect 57099 652900 57165 652901
rect 57099 652836 57100 652900
rect 57164 652836 57165 652900
rect 57099 652835 57165 652836
rect 57102 42533 57162 652835
rect 57651 147796 57717 147797
rect 57651 147732 57652 147796
rect 57716 147732 57717 147796
rect 57651 147731 57717 147732
rect 57099 42532 57165 42533
rect 57099 42468 57100 42532
rect 57164 42468 57165 42532
rect 57099 42467 57165 42468
rect 56363 41308 56429 41309
rect 56363 41244 56364 41308
rect 56428 41244 56429 41308
rect 56363 41243 56429 41244
rect 56179 6628 56245 6629
rect 56179 6564 56180 6628
rect 56244 6564 56245 6628
rect 56179 6563 56245 6564
rect 57654 6493 57714 147731
rect 57838 41173 57898 700435
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 267005 73404 289898
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 267005 91404 271898
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 267005 109404 289898
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 267005 127404 271898
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 267005 145404 289898
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 267005 163404 271898
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 267005 181404 289898
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 267005 199404 271898
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 267005 217404 289898
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 267005 235404 271898
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 241467 267340 241533 267341
rect 241467 267276 241468 267340
rect 241532 267276 241533 267340
rect 241467 267275 241533 267276
rect 244595 267340 244661 267341
rect 244595 267276 244596 267340
rect 244660 267276 244661 267340
rect 244595 267275 244661 267276
rect 241470 267018 241530 267275
rect 244598 267018 244658 267275
rect 252804 267005 253404 289898
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 285627 700364 285693 700365
rect 285627 700300 285628 700364
rect 285692 700300 285693 700364
rect 285627 700299 285693 700300
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 267005 271404 271898
rect 280475 269652 280541 269653
rect 280475 269588 280476 269652
rect 280540 269588 280541 269652
rect 280475 269587 280541 269588
rect 278819 269516 278885 269517
rect 278819 269452 278820 269516
rect 278884 269452 278885 269516
rect 278819 269451 278885 269452
rect 278635 267340 278701 267341
rect 278635 267276 278636 267340
rect 278700 267276 278701 267340
rect 278635 267275 278701 267276
rect 64643 266524 64709 266525
rect 64643 266460 64644 266524
rect 64708 266460 64709 266524
rect 64643 266459 64709 266460
rect 64459 264348 64525 264349
rect 64459 264284 64460 264348
rect 64524 264284 64525 264348
rect 64459 264283 64525 264284
rect 63355 263668 63421 263669
rect 63355 263604 63356 263668
rect 63420 263604 63421 263668
rect 63355 263603 63421 263604
rect 60779 247348 60845 247349
rect 60779 247284 60780 247348
rect 60844 247284 60845 247348
rect 60779 247283 60845 247284
rect 59675 228308 59741 228309
rect 59675 228244 59676 228308
rect 59740 228244 59741 228308
rect 59675 228243 59741 228244
rect 59123 200564 59189 200565
rect 59123 200500 59124 200564
rect 59188 200500 59189 200564
rect 59123 200499 59189 200500
rect 58755 171188 58821 171189
rect 58755 171124 58756 171188
rect 58820 171124 58821 171188
rect 58755 171123 58821 171124
rect 58571 144804 58637 144805
rect 58571 144740 58572 144804
rect 58636 144740 58637 144804
rect 58571 144739 58637 144740
rect 57835 41172 57901 41173
rect 57835 41108 57836 41172
rect 57900 41108 57901 41172
rect 57835 41107 57901 41108
rect 58574 15877 58634 144739
rect 58758 24173 58818 171123
rect 58939 161124 59005 161125
rect 58939 161060 58940 161124
rect 59004 161060 59005 161124
rect 58939 161059 59005 161060
rect 58755 24172 58821 24173
rect 58755 24108 58756 24172
rect 58820 24108 58821 24172
rect 58755 24107 58821 24108
rect 58571 15876 58637 15877
rect 58571 15812 58572 15876
rect 58636 15812 58637 15876
rect 58571 15811 58637 15812
rect 57651 6492 57717 6493
rect 57651 6428 57652 6492
rect 57716 6428 57717 6492
rect 57651 6427 57717 6428
rect 58942 4861 59002 161059
rect 59126 32469 59186 200499
rect 59307 137732 59373 137733
rect 59307 137668 59308 137732
rect 59372 137668 59373 137732
rect 59307 137667 59373 137668
rect 59123 32468 59189 32469
rect 59123 32404 59124 32468
rect 59188 32404 59189 32468
rect 59123 32403 59189 32404
rect 59310 25533 59370 137667
rect 59678 68458 59738 228243
rect 60595 210628 60661 210629
rect 60595 210564 60596 210628
rect 60660 210564 60661 210628
rect 60595 210563 60661 210564
rect 60043 109716 60109 109717
rect 60043 109652 60044 109716
rect 60108 109652 60109 109716
rect 60043 109651 60109 109652
rect 60046 69138 60106 109651
rect 60411 75852 60477 75853
rect 60411 75788 60412 75852
rect 60476 75788 60477 75852
rect 60411 75787 60477 75788
rect 60043 61572 60109 61573
rect 60043 61508 60044 61572
rect 60108 61508 60109 61572
rect 60043 61507 60109 61508
rect 60046 29613 60106 61507
rect 60414 32605 60474 75787
rect 60598 33829 60658 210563
rect 60595 33828 60661 33829
rect 60595 33764 60596 33828
rect 60660 33764 60661 33828
rect 60595 33763 60661 33764
rect 60411 32604 60477 32605
rect 60411 32540 60412 32604
rect 60476 32540 60477 32604
rect 60411 32539 60477 32540
rect 60782 29749 60842 247283
rect 60966 194309 61026 249102
rect 60963 194308 61029 194309
rect 60963 194244 60964 194308
rect 61028 194244 61029 194308
rect 60963 194243 61029 194244
rect 61334 180709 61394 251142
rect 61702 208045 61762 248422
rect 62619 243812 62685 243813
rect 62619 243748 62620 243812
rect 62684 243748 62685 243812
rect 62619 243747 62685 243748
rect 62622 234970 62682 243747
rect 63358 240274 63418 263603
rect 63358 240214 63602 240274
rect 63542 239730 63602 240214
rect 63358 239670 63602 239730
rect 63358 239050 63418 239670
rect 62438 234910 62682 234970
rect 63174 238990 63418 239050
rect 62438 224770 62498 234910
rect 62438 224710 62682 224770
rect 61883 208316 61949 208317
rect 61883 208252 61884 208316
rect 61948 208252 61949 208316
rect 61883 208251 61949 208252
rect 61699 208044 61765 208045
rect 61699 207980 61700 208044
rect 61764 207980 61765 208044
rect 61699 207979 61765 207980
rect 61699 193356 61765 193357
rect 61699 193292 61700 193356
rect 61764 193292 61765 193356
rect 61699 193291 61765 193292
rect 61331 180708 61397 180709
rect 61331 180644 61332 180708
rect 61396 180644 61397 180708
rect 61331 180643 61397 180644
rect 61147 81564 61213 81565
rect 61147 81500 61148 81564
rect 61212 81500 61213 81564
rect 61147 81499 61213 81500
rect 61150 72538 61210 81499
rect 61515 73132 61581 73133
rect 61515 73068 61516 73132
rect 61580 73068 61581 73132
rect 61515 73067 61581 73068
rect 61518 36549 61578 73067
rect 61515 36548 61581 36549
rect 61515 36484 61516 36548
rect 61580 36484 61581 36548
rect 61515 36483 61581 36484
rect 61702 35189 61762 193291
rect 61699 35188 61765 35189
rect 61699 35124 61700 35188
rect 61764 35124 61765 35188
rect 61699 35123 61765 35124
rect 60779 29748 60845 29749
rect 60779 29684 60780 29748
rect 60844 29684 60845 29748
rect 60779 29683 60845 29684
rect 60043 29612 60109 29613
rect 60043 29548 60044 29612
rect 60108 29548 60109 29612
rect 60043 29547 60109 29548
rect 59307 25532 59373 25533
rect 59307 25468 59308 25532
rect 59372 25468 59373 25532
rect 59307 25467 59373 25468
rect 61886 21317 61946 208251
rect 62622 205869 62682 224710
rect 63174 222050 63234 238990
rect 62990 221990 63234 222050
rect 62990 220690 63050 221990
rect 62806 220630 63050 220690
rect 62806 212258 62866 220630
rect 62806 212198 63602 212258
rect 63542 211170 63602 212198
rect 63358 211110 63602 211170
rect 62619 205868 62685 205869
rect 62619 205804 62620 205868
rect 62684 205804 62685 205868
rect 62619 205803 62685 205804
rect 63358 201650 63418 211110
rect 63174 201590 63418 201650
rect 62619 201516 62685 201517
rect 62619 201452 62620 201516
rect 62684 201452 62685 201516
rect 62619 201451 62685 201452
rect 62622 183837 62682 201451
rect 63174 196210 63234 201590
rect 63174 196150 63602 196210
rect 63542 190770 63602 196150
rect 63542 190710 64338 190770
rect 62619 183836 62685 183837
rect 62619 183772 62620 183836
rect 62684 183772 62685 183836
rect 62619 183771 62685 183772
rect 62435 183700 62501 183701
rect 62435 183636 62436 183700
rect 62500 183636 62501 183700
rect 62435 183635 62501 183636
rect 62438 154597 62498 183635
rect 64278 183290 64338 190710
rect 64094 183230 64338 183290
rect 64094 182610 64154 183230
rect 63910 182550 64154 182610
rect 63910 177170 63970 182550
rect 63358 177110 63970 177170
rect 63358 173770 63418 177110
rect 63358 173710 63602 173770
rect 62619 157180 62685 157181
rect 62619 157116 62620 157180
rect 62684 157116 62685 157180
rect 62619 157115 62685 157116
rect 62067 154596 62133 154597
rect 62067 154532 62068 154596
rect 62132 154532 62133 154596
rect 62067 154531 62133 154532
rect 62435 154596 62501 154597
rect 62435 154532 62436 154596
rect 62500 154532 62501 154596
rect 62435 154531 62501 154532
rect 62070 143717 62130 154531
rect 62622 143850 62682 157115
rect 63542 154050 63602 173710
rect 63174 153990 63602 154050
rect 63174 149290 63234 153990
rect 63174 149230 63602 149290
rect 62622 143790 63050 143850
rect 62067 143716 62133 143717
rect 62067 143652 62068 143716
rect 62132 143652 62133 143716
rect 62067 143651 62133 143652
rect 62619 143580 62685 143581
rect 62619 143516 62620 143580
rect 62684 143516 62685 143580
rect 62619 143515 62685 143516
rect 62622 137050 62682 143515
rect 62254 136990 62682 137050
rect 62254 128213 62314 136990
rect 62990 135146 63050 143790
rect 62622 135086 63050 135146
rect 62251 128212 62317 128213
rect 62251 128148 62252 128212
rect 62316 128148 62317 128212
rect 62251 128147 62317 128148
rect 62622 128077 62682 135086
rect 63542 128210 63602 149230
rect 63358 128150 63602 128210
rect 62251 128076 62317 128077
rect 62251 128012 62252 128076
rect 62316 128012 62317 128076
rect 62251 128011 62317 128012
rect 62619 128076 62685 128077
rect 62619 128012 62620 128076
rect 62684 128012 62685 128076
rect 62619 128011 62685 128012
rect 62254 117333 62314 128011
rect 63358 125490 63418 128150
rect 63358 125430 63786 125490
rect 62251 117332 62317 117333
rect 62251 117268 62252 117332
rect 62316 117268 62317 117332
rect 62251 117267 62317 117268
rect 62619 117332 62685 117333
rect 62619 117268 62620 117332
rect 62684 117330 62685 117332
rect 62684 117270 63234 117330
rect 62684 117268 62685 117270
rect 62619 117267 62685 117268
rect 62435 115972 62501 115973
rect 62435 115908 62436 115972
rect 62500 115970 62501 115972
rect 63174 115970 63234 117270
rect 63726 115970 63786 125430
rect 62500 115910 62682 115970
rect 62500 115908 62501 115910
rect 62435 115907 62501 115908
rect 62622 111485 62682 115910
rect 62806 115910 63234 115970
rect 63358 115910 63786 115970
rect 62619 111484 62685 111485
rect 62619 111420 62620 111484
rect 62684 111420 62685 111484
rect 62619 111419 62685 111420
rect 62806 110530 62866 115910
rect 63358 110530 63418 115910
rect 62438 110470 62866 110530
rect 62990 110470 63418 110530
rect 62438 93530 62498 110470
rect 62619 106316 62685 106317
rect 62619 106252 62620 106316
rect 62684 106252 62685 106316
rect 62619 106251 62685 106252
rect 62622 106045 62682 106251
rect 62619 106044 62685 106045
rect 62619 105980 62620 106044
rect 62684 105980 62685 106044
rect 62619 105979 62685 105980
rect 62990 102370 63050 110470
rect 62990 102310 63234 102370
rect 63174 101010 63234 102310
rect 63174 100950 63602 101010
rect 62619 98292 62685 98293
rect 62619 98228 62620 98292
rect 62684 98228 62685 98292
rect 62619 98227 62685 98228
rect 62622 93805 62682 98227
rect 63542 96930 63602 100950
rect 63174 96870 63602 96930
rect 62619 93804 62685 93805
rect 62619 93740 62620 93804
rect 62684 93740 62685 93804
rect 63174 93802 63234 96870
rect 63174 93742 63786 93802
rect 62619 93739 62685 93740
rect 62438 93470 63234 93530
rect 62619 88636 62685 88637
rect 62619 88572 62620 88636
rect 62684 88572 62685 88636
rect 62619 88571 62685 88572
rect 62622 83330 62682 88571
rect 63174 88090 63234 93470
rect 62438 83270 62682 83330
rect 62806 88030 63234 88090
rect 62438 79250 62498 83270
rect 62619 79932 62685 79933
rect 62619 79868 62620 79932
rect 62684 79930 62685 79932
rect 62806 79930 62866 88030
rect 63726 87410 63786 93742
rect 63358 87350 63786 87410
rect 63358 84010 63418 87350
rect 63358 83950 63602 84010
rect 62684 79870 62866 79930
rect 62684 79868 62685 79870
rect 62619 79867 62685 79868
rect 62438 79190 62682 79250
rect 62622 70549 62682 79190
rect 62619 70548 62685 70549
rect 62619 70484 62620 70548
rect 62684 70484 62685 70548
rect 62619 70483 62685 70484
rect 63542 70410 63602 83950
rect 63358 70350 63602 70410
rect 62619 67828 62685 67829
rect 62619 67764 62620 67828
rect 62684 67764 62685 67828
rect 62619 67763 62685 67764
rect 62622 65650 62682 67763
rect 62622 65590 62866 65650
rect 62806 60890 62866 65590
rect 62806 60830 63234 60890
rect 62619 60756 62685 60757
rect 62619 60692 62620 60756
rect 62684 60692 62685 60756
rect 62619 60691 62685 60692
rect 62622 52461 62682 60691
rect 63174 54770 63234 60830
rect 62806 54710 63234 54770
rect 62067 52460 62133 52461
rect 62067 52396 62068 52460
rect 62132 52396 62133 52460
rect 62067 52395 62133 52396
rect 62619 52460 62685 52461
rect 62619 52396 62620 52460
rect 62684 52396 62685 52460
rect 62619 52395 62685 52396
rect 62070 43757 62130 52395
rect 62251 48244 62317 48245
rect 62251 48180 62252 48244
rect 62316 48180 62317 48244
rect 62251 48179 62317 48180
rect 62254 43893 62314 48179
rect 62806 47970 62866 54710
rect 63358 48650 63418 70350
rect 63726 52050 63786 68902
rect 64094 64970 64154 68222
rect 64094 64910 64338 64970
rect 64278 52050 64338 64910
rect 63542 51990 63786 52050
rect 63910 51990 64338 52050
rect 63542 49330 63602 51990
rect 63542 49270 63786 49330
rect 63358 48590 63602 48650
rect 62438 47910 62866 47970
rect 62251 43892 62317 43893
rect 62251 43828 62252 43892
rect 62316 43828 62317 43892
rect 62251 43827 62317 43828
rect 62067 43756 62133 43757
rect 62067 43692 62068 43756
rect 62132 43692 62133 43756
rect 62067 43691 62133 43692
rect 62438 37909 62498 47910
rect 63542 43893 63602 48590
rect 62987 43892 63053 43893
rect 62987 43828 62988 43892
rect 63052 43828 63053 43892
rect 62987 43827 63053 43828
rect 63539 43892 63605 43893
rect 63539 43828 63540 43892
rect 63604 43828 63605 43892
rect 63539 43827 63605 43828
rect 62803 43756 62869 43757
rect 62803 43692 62804 43756
rect 62868 43692 62869 43756
rect 62803 43691 62869 43692
rect 62806 41170 62866 43691
rect 62622 41110 62866 41170
rect 62435 37908 62501 37909
rect 62435 37844 62436 37908
rect 62500 37844 62501 37908
rect 62435 37843 62501 37844
rect 62622 30973 62682 41110
rect 62619 30972 62685 30973
rect 62619 30908 62620 30972
rect 62684 30908 62685 30972
rect 62619 30907 62685 30908
rect 62990 25669 63050 43827
rect 62987 25668 63053 25669
rect 62987 25604 62988 25668
rect 63052 25604 63053 25668
rect 62987 25603 63053 25604
rect 61883 21316 61949 21317
rect 61883 21252 61884 21316
rect 61948 21252 61949 21316
rect 61883 21251 61949 21252
rect 58939 4860 59005 4861
rect 58939 4796 58940 4860
rect 59004 4796 59005 4860
rect 58939 4795 59005 4796
rect 63726 3229 63786 49270
rect 63910 41170 63970 51990
rect 63910 41110 64154 41170
rect 64094 31925 64154 41110
rect 64091 31924 64157 31925
rect 64091 31860 64092 31924
rect 64156 31860 64157 31924
rect 64091 31859 64157 31860
rect 64275 31788 64341 31789
rect 64275 31724 64276 31788
rect 64340 31724 64341 31788
rect 64275 31723 64341 31724
rect 64278 19413 64338 31723
rect 64462 28253 64522 264283
rect 64459 28252 64525 28253
rect 64459 28188 64460 28252
rect 64524 28188 64525 28252
rect 64459 28187 64525 28188
rect 64275 19412 64341 19413
rect 64275 19348 64276 19412
rect 64340 19348 64341 19412
rect 64275 19347 64341 19348
rect 64275 19140 64341 19141
rect 64275 19076 64276 19140
rect 64340 19076 64341 19140
rect 64275 19075 64341 19076
rect 64278 11930 64338 19075
rect 63910 11870 64338 11930
rect 63910 3773 63970 11870
rect 63907 3772 63973 3773
rect 63907 3708 63908 3772
rect 63972 3708 63973 3772
rect 63907 3707 63973 3708
rect 64646 3637 64706 266459
rect 231902 266253 231962 266782
rect 231899 266252 231965 266253
rect 231899 266188 231900 266252
rect 231964 266188 231965 266252
rect 231899 266187 231965 266188
rect 155907 264348 155973 264349
rect 155907 264284 155908 264348
rect 155972 264284 155973 264348
rect 155907 264283 155973 264284
rect 201723 264348 201789 264349
rect 201723 264284 201724 264348
rect 201788 264284 201789 264348
rect 201723 264283 201789 264284
rect 224907 264348 224973 264349
rect 224907 264284 224908 264348
rect 224972 264284 224973 264348
rect 224907 264283 224973 264284
rect 259131 264348 259197 264349
rect 259131 264284 259132 264348
rect 259196 264284 259197 264348
rect 259131 264283 259197 264284
rect 155910 263669 155970 264283
rect 155907 263668 155973 263669
rect 155907 263604 155908 263668
rect 155972 263604 155973 263668
rect 155907 263603 155973 263604
rect 201726 262938 201786 264283
rect 224910 264077 224970 264283
rect 224907 264076 224973 264077
rect 224907 264012 224908 264076
rect 224972 264012 224973 264076
rect 224907 264011 224973 264012
rect 259134 263805 259194 264283
rect 259131 263804 259197 263805
rect 259131 263740 259132 263804
rect 259196 263740 259197 263804
rect 259131 263739 259197 263740
rect 278638 263533 278698 267275
rect 278635 263532 278701 263533
rect 278635 263468 278636 263532
rect 278700 263468 278701 263532
rect 278635 263467 278701 263468
rect 65379 43892 65445 43893
rect 65379 43828 65380 43892
rect 65444 43828 65445 43892
rect 65379 43827 65445 43828
rect 65382 6901 65442 43827
rect 276982 42261 277042 44422
rect 277163 43892 277229 43893
rect 277163 43828 277164 43892
rect 277228 43828 277229 43892
rect 277163 43827 277229 43828
rect 276979 42260 277045 42261
rect 276979 42196 276980 42260
rect 277044 42196 277045 42260
rect 276979 42195 277045 42196
rect 72804 38454 73404 41200
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 65379 6900 65445 6901
rect 65379 6836 65380 6900
rect 65444 6836 65445 6900
rect 65379 6835 65445 6836
rect 64643 3636 64709 3637
rect 64643 3572 64644 3636
rect 64708 3572 64709 3636
rect 64643 3571 64709 3572
rect 63723 3228 63789 3229
rect 63723 3164 63724 3228
rect 63788 3164 63789 3228
rect 63723 3163 63789 3164
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 90804 20454 91404 41200
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 108804 38454 109404 41200
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 126804 20454 127404 41200
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 144804 38454 145404 41200
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 162804 20454 163404 41200
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 180804 38454 181404 41200
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 198804 20454 199404 41200
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 216804 38454 217404 41200
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 234804 20454 235404 41200
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 252804 38454 253404 41200
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 270804 20454 271404 41200
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 277166 6901 277226 43827
rect 278822 39405 278882 269451
rect 280107 267612 280173 267613
rect 280107 267548 280108 267612
rect 280172 267548 280173 267612
rect 280107 267547 280173 267548
rect 280110 267018 280170 267547
rect 279371 264348 279437 264349
rect 279371 264284 279372 264348
rect 279436 264284 279437 264348
rect 279371 264283 279437 264284
rect 278819 39404 278885 39405
rect 278819 39340 278820 39404
rect 278884 39340 278885 39404
rect 278819 39339 278885 39340
rect 277163 6900 277229 6901
rect 277163 6836 277164 6900
rect 277228 6836 277229 6900
rect 277163 6835 277229 6836
rect 279374 3229 279434 264283
rect 279742 3637 279802 60742
rect 280478 39269 280538 269587
rect 282499 269380 282565 269381
rect 282499 269316 282500 269380
rect 282564 269316 282565 269380
rect 282499 269315 282565 269316
rect 281763 268020 281829 268021
rect 281763 267956 281764 268020
rect 281828 267956 281829 268020
rect 281763 267955 281829 267956
rect 280659 265708 280725 265709
rect 280659 265644 280660 265708
rect 280724 265644 280725 265708
rect 280659 265643 280725 265644
rect 280475 39268 280541 39269
rect 280475 39204 280476 39268
rect 280540 39204 280541 39268
rect 280475 39203 280541 39204
rect 280662 3637 280722 265643
rect 280843 265028 280909 265029
rect 280843 264964 280844 265028
rect 280908 264964 280909 265028
rect 280843 264963 280909 264964
rect 280846 3773 280906 264963
rect 281027 264076 281093 264077
rect 281027 264012 281028 264076
rect 281092 264012 281093 264076
rect 281027 264011 281093 264012
rect 281030 4045 281090 264011
rect 281579 214436 281645 214437
rect 281579 214372 281580 214436
rect 281644 214372 281645 214436
rect 281579 214371 281645 214372
rect 281582 79250 281642 214371
rect 281398 79190 281642 79250
rect 281398 77978 281458 79190
rect 281766 43485 281826 267955
rect 282131 248372 282132 248422
rect 282196 248372 282197 248422
rect 282131 248371 282197 248372
rect 282131 126988 282197 126989
rect 282131 126924 282132 126988
rect 282196 126924 282197 126988
rect 282131 126923 282197 126924
rect 281947 52460 282013 52461
rect 281947 52396 281948 52460
rect 282012 52396 282013 52460
rect 281947 52395 282013 52396
rect 281763 43484 281829 43485
rect 281763 43420 281764 43484
rect 281828 43420 281829 43484
rect 281763 43419 281829 43420
rect 281950 40901 282010 52395
rect 281947 40900 282013 40901
rect 281947 40836 281948 40900
rect 282012 40836 282013 40900
rect 281947 40835 282013 40836
rect 281027 4044 281093 4045
rect 281027 3980 281028 4044
rect 281092 3980 281093 4044
rect 281027 3979 281093 3980
rect 282134 3909 282194 126923
rect 282502 44658 282562 269315
rect 282867 256052 282933 256053
rect 282867 255988 282868 256052
rect 282932 255988 282933 256052
rect 282867 255987 282933 255988
rect 282870 16013 282930 255987
rect 283235 244220 283301 244221
rect 283235 244156 283236 244220
rect 283300 244156 283301 244220
rect 283235 244155 283301 244156
rect 283238 241501 283298 244155
rect 283235 241500 283301 241501
rect 283235 241436 283236 241500
rect 283300 241436 283301 241500
rect 283235 241435 283301 241436
rect 283422 221509 283482 251142
rect 283603 248436 283669 248437
rect 283603 248372 283604 248436
rect 283668 248372 283669 248436
rect 283603 248371 283669 248372
rect 283606 244221 283666 248371
rect 283603 244220 283669 244221
rect 283603 244156 283604 244220
rect 283668 244156 283669 244220
rect 283603 244155 283669 244156
rect 283974 234837 284034 250462
rect 283971 234836 284037 234837
rect 283971 234772 283972 234836
rect 284036 234772 284037 234836
rect 283971 234771 284037 234772
rect 283787 232116 283853 232117
rect 283787 232052 283788 232116
rect 283852 232052 283853 232116
rect 283787 232051 283853 232052
rect 283603 231980 283669 231981
rect 283603 231916 283604 231980
rect 283668 231916 283669 231980
rect 283603 231915 283669 231916
rect 283419 221508 283485 221509
rect 283419 221444 283420 221508
rect 283484 221444 283485 221508
rect 283419 221443 283485 221444
rect 283419 221236 283485 221237
rect 283419 221172 283420 221236
rect 283484 221172 283485 221236
rect 283419 221171 283485 221172
rect 283235 220148 283301 220149
rect 283235 220084 283236 220148
rect 283300 220084 283301 220148
rect 283235 220083 283301 220084
rect 283051 209676 283117 209677
rect 283051 209612 283052 209676
rect 283116 209612 283117 209676
rect 283051 209611 283117 209612
rect 283054 41037 283114 209611
rect 283238 206277 283298 220083
rect 283422 209269 283482 221171
rect 283606 220149 283666 231915
rect 283603 220148 283669 220149
rect 283603 220084 283604 220148
rect 283668 220084 283669 220148
rect 283603 220083 283669 220084
rect 283790 220010 283850 232051
rect 283606 219950 283850 220010
rect 283606 209405 283666 219950
rect 283603 209404 283669 209405
rect 283603 209340 283604 209404
rect 283668 209340 283669 209404
rect 283603 209339 283669 209340
rect 283419 209268 283485 209269
rect 283419 209204 283420 209268
rect 283484 209204 283485 209268
rect 283419 209203 283485 209204
rect 283419 208996 283485 208997
rect 283419 208932 283420 208996
rect 283484 208932 283485 208996
rect 283419 208931 283485 208932
rect 283235 206276 283301 206277
rect 283235 206212 283236 206276
rect 283300 206212 283301 206276
rect 283235 206211 283301 206212
rect 283235 180436 283301 180437
rect 283235 180372 283236 180436
rect 283300 180372 283301 180436
rect 283235 180371 283301 180372
rect 283238 174589 283298 180371
rect 283235 174588 283301 174589
rect 283235 174524 283236 174588
rect 283300 174524 283301 174588
rect 283235 174523 283301 174524
rect 283422 168197 283482 208931
rect 283971 206276 284037 206277
rect 283971 206212 283972 206276
rect 284036 206212 284037 206276
rect 283971 206211 284037 206212
rect 283974 192541 284034 206211
rect 283971 192540 284037 192541
rect 283971 192476 283972 192540
rect 284036 192476 284037 192540
rect 283971 192475 284037 192476
rect 283787 174588 283853 174589
rect 283787 174524 283788 174588
rect 283852 174524 283853 174588
rect 283787 174523 283853 174524
rect 283419 168196 283485 168197
rect 283419 168132 283420 168196
rect 283484 168132 283485 168196
rect 283419 168131 283485 168132
rect 283790 162485 283850 174523
rect 283787 162484 283853 162485
rect 283787 162420 283788 162484
rect 283852 162420 283853 162484
rect 283787 162419 283853 162420
rect 283422 72453 283482 72982
rect 283419 72452 283485 72453
rect 283419 72388 283420 72452
rect 283484 72388 283485 72452
rect 283419 72387 283485 72388
rect 283235 52596 283301 52597
rect 283235 52532 283236 52596
rect 283300 52532 283301 52596
rect 283235 52531 283301 52532
rect 283051 41036 283117 41037
rect 283051 40972 283052 41036
rect 283116 40972 283117 41036
rect 283051 40971 283117 40972
rect 283238 29885 283298 52531
rect 283235 29884 283301 29885
rect 283235 29820 283236 29884
rect 283300 29820 283301 29884
rect 283235 29819 283301 29820
rect 282867 16012 282933 16013
rect 282867 15948 282868 16012
rect 282932 15948 282933 16012
rect 282867 15947 282933 15948
rect 284342 6085 284402 262702
rect 285630 41173 285690 700299
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 286179 556204 286245 556205
rect 286179 556140 286180 556204
rect 286244 556140 286245 556204
rect 286179 556139 286245 556140
rect 286182 42669 286242 556139
rect 288804 542454 289404 577898
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 299611 569940 299677 569941
rect 299611 569876 299612 569940
rect 299676 569876 299677 569940
rect 299611 569875 299677 569876
rect 299614 560421 299674 569875
rect 306804 560454 307404 595898
rect 299611 560420 299677 560421
rect 299611 560356 299612 560420
rect 299676 560356 299677 560420
rect 299611 560355 299677 560356
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 299427 556476 299493 556477
rect 299427 556412 299428 556476
rect 299492 556412 299493 556476
rect 299427 556411 299493 556412
rect 299430 556205 299490 556411
rect 299427 556204 299493 556205
rect 299427 556140 299428 556204
rect 299492 556140 299493 556204
rect 299427 556139 299493 556140
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 299611 273324 299677 273325
rect 299611 273260 299612 273324
rect 299676 273260 299677 273324
rect 299611 273259 299677 273260
rect 299614 270605 299674 273259
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 299611 270604 299677 270605
rect 299611 270540 299612 270604
rect 299676 270540 299677 270604
rect 299611 270539 299677 270540
rect 294643 267612 294709 267613
rect 294643 267548 294644 267612
rect 294708 267548 294709 267612
rect 294643 267547 294709 267548
rect 294646 267018 294706 267547
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 306804 236454 307404 271898
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 308995 266932 309061 266933
rect 308995 266868 308996 266932
rect 309060 266868 309061 266932
rect 308995 266867 309061 266868
rect 308998 266338 309058 266867
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 297958 76533 298018 77062
rect 297955 76532 298021 76533
rect 297955 76468 297956 76532
rect 298020 76468 298021 76532
rect 297955 76467 298021 76468
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 286179 42668 286245 42669
rect 286179 42604 286180 42668
rect 286244 42604 286245 42668
rect 286179 42603 286245 42604
rect 285627 41172 285693 41173
rect 285627 41108 285628 41172
rect 285692 41108 285693 41172
rect 285627 41107 285693 41108
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 284339 6084 284405 6085
rect 284339 6020 284340 6084
rect 284404 6020 284405 6084
rect 284339 6019 284405 6020
rect 282131 3908 282197 3909
rect 282131 3844 282132 3908
rect 282196 3844 282197 3908
rect 282131 3843 282197 3844
rect 280843 3772 280909 3773
rect 280843 3708 280844 3772
rect 280908 3708 280909 3772
rect 280843 3707 280909 3708
rect 279739 3636 279805 3637
rect 279739 3572 279740 3636
rect 279804 3572 279805 3636
rect 279739 3571 279805 3572
rect 280659 3636 280725 3637
rect 280659 3572 280660 3636
rect 280724 3572 280725 3636
rect 280659 3571 280725 3572
rect 279371 3228 279437 3229
rect 279371 3164 279372 3228
rect 279436 3164 279437 3228
rect 279371 3163 279437 3164
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 306804 56454 307404 91898
rect 324804 254454 325404 289898
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 328315 266932 328381 266933
rect 328315 266868 328316 266932
rect 328380 266868 328381 266932
rect 328315 266867 328381 266868
rect 328318 266338 328378 266867
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 318566 71773 318626 72302
rect 318563 71772 318629 71773
rect 318563 71708 318564 71772
rect 318628 71708 318629 71772
rect 318563 71707 318629 71708
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 324804 38454 325404 73898
rect 342804 236454 343404 271898
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 347635 266932 347701 266933
rect 347635 266868 347636 266932
rect 347700 266868 347701 266932
rect 347635 266867 347701 266868
rect 347638 266338 347698 266867
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 337886 71773 337946 72302
rect 337883 71772 337949 71773
rect 337883 71708 337884 71772
rect 337948 71708 337949 71772
rect 337883 71707 337949 71708
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 342804 56454 343404 91898
rect 360804 254454 361404 289898
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 366955 266932 367021 266933
rect 366955 266868 366956 266932
rect 367020 266868 367021 266932
rect 366955 266867 367021 266868
rect 366958 266338 367018 266867
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 357206 75853 357266 76382
rect 357203 75852 357269 75853
rect 357203 75788 357204 75852
rect 357268 75788 357269 75852
rect 357203 75787 357269 75788
rect 360804 74454 361404 109898
rect 378804 236454 379404 271898
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 386275 266932 386341 266933
rect 386275 266868 386276 266932
rect 386340 266868 386341 266932
rect 386275 266867 386341 266868
rect 386278 266338 386338 266867
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 357206 71773 357266 72302
rect 357203 71772 357269 71773
rect 357203 71708 357204 71772
rect 357268 71708 357269 71772
rect 357203 71707 357269 71708
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 360804 38454 361404 73898
rect 376526 71773 376586 72302
rect 376523 71772 376589 71773
rect 376523 71708 376524 71772
rect 376588 71708 376589 71772
rect 376523 71707 376589 71708
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 378804 56454 379404 91898
rect 396804 254454 397404 289898
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 405595 266932 405661 266933
rect 405595 266868 405596 266932
rect 405660 266868 405661 266932
rect 405595 266867 405661 266868
rect 405598 266338 405658 266867
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 386278 72453 386338 72982
rect 386275 72452 386341 72453
rect 386275 72388 386276 72452
rect 386340 72388 386341 72452
rect 386275 72387 386341 72388
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 396804 38454 397404 73898
rect 414804 236454 415404 271898
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 434667 556476 434733 556477
rect 434667 556412 434668 556476
rect 434732 556412 434733 556476
rect 434667 556411 434733 556412
rect 434670 555933 434730 556411
rect 434667 555932 434733 555933
rect 434667 555868 434668 555932
rect 434732 555868 434733 555932
rect 434667 555867 434733 555868
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 424915 266932 424981 266933
rect 424915 266868 424916 266932
rect 424980 266868 424981 266932
rect 424915 266867 424981 266868
rect 424918 266338 424978 266867
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 405782 69818 405842 71622
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 414804 56454 415404 91898
rect 432804 254454 433404 289898
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 444235 266932 444301 266933
rect 444235 266868 444236 266932
rect 444300 266868 444301 266932
rect 444235 266867 444301 266868
rect 444238 266338 444298 266867
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 424915 72452 424981 72453
rect 424915 72388 424916 72452
rect 424980 72388 424981 72452
rect 424915 72387 424981 72388
rect 424918 71858 424978 72387
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 432804 38454 433404 73898
rect 450804 236454 451404 271898
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 463555 266932 463621 266933
rect 463555 266868 463556 266932
rect 463620 266868 463621 266932
rect 463555 266867 463621 266868
rect 463558 266338 463618 266867
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 450804 56454 451404 91898
rect 468804 254454 469404 289898
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 482875 266932 482941 266933
rect 482875 266868 482876 266932
rect 482940 266868 482941 266932
rect 482875 266867 482941 266868
rect 482878 266338 482938 266867
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 468804 38454 469404 73898
rect 486804 236454 487404 271898
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 502195 266932 502261 266933
rect 502195 266868 502196 266932
rect 502260 266868 502261 266932
rect 502195 266867 502261 266868
rect 502198 266338 502258 266867
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 486804 56454 487404 91898
rect 504804 254454 505404 289898
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 521515 266932 521581 266933
rect 521515 266868 521516 266932
rect 521580 266868 521581 266932
rect 521515 266867 521581 266868
rect 521518 266338 521578 266867
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 500723 77212 500789 77213
rect 500723 77148 500724 77212
rect 500788 77148 500789 77212
rect 500723 77147 500789 77148
rect 500726 76618 500786 77147
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 504804 38454 505404 73898
rect 522804 236454 523404 271898
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 533846 266933 533906 267462
rect 533843 266932 533909 266933
rect 533843 266868 533844 266932
rect 533908 266868 533909 266932
rect 533843 266867 533909 266868
rect 536787 266932 536853 266933
rect 536787 266868 536788 266932
rect 536852 266868 536853 266932
rect 536787 266867 536853 266868
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 536790 3501 536850 266867
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 542675 80068 542741 80069
rect 542675 80004 542676 80068
rect 542740 80004 542741 80068
rect 542675 80003 542741 80004
rect 542678 77349 542738 80003
rect 542675 77348 542741 77349
rect 542675 77284 542676 77348
rect 542740 77284 542741 77348
rect 542675 77283 542741 77284
rect 542491 77212 542557 77213
rect 542491 77148 542492 77212
rect 542556 77148 542557 77212
rect 542491 77147 542557 77148
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 542494 67693 542554 77147
rect 542491 67692 542557 67693
rect 542491 67628 542492 67692
rect 542556 67628 542557 67692
rect 542491 67627 542557 67628
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 536787 3500 536853 3501
rect 536787 3436 536788 3500
rect 536852 3436 536853 3500
rect 536787 3435 536853 3436
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 576804 704838 577404 705800
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 580763 217020 580829 217021
rect 580763 216956 580764 217020
rect 580828 216956 580829 217020
rect 580763 216955 580829 216956
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 580395 111484 580461 111485
rect 580395 111420 580396 111484
rect 580460 111420 580461 111484
rect 580395 111419 580461 111420
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 580398 73218 580458 111419
rect 580766 76618 580826 216955
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 587200 -2226 587800 706162
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 588140 -3166 588740 707102
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 589080 -4106 589680 708042
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 590020 -5046 590620 708982
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 590960 -5986 591560 709922
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 591900 -6926 592500 710862
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 3286 79102 3522 79338
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 22606 79252 22842 79338
rect 22606 79188 22692 79252
rect 22692 79188 22756 79252
rect 22756 79188 22842 79252
rect 22606 79102 22842 79188
rect 28862 79252 29098 79338
rect 28862 79188 28948 79252
rect 28948 79188 29012 79252
rect 29012 79188 29098 79252
rect 28862 79102 29098 79188
rect 19478 77742 19714 77978
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 41926 79252 42162 79338
rect 41926 79188 42012 79252
rect 42012 79188 42076 79252
rect 42076 79188 42162 79252
rect 41926 79102 42162 79188
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 107430 266932 107666 267018
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 107430 266868 107516 266932
rect 107516 266868 107580 266932
rect 107580 266868 107666 266932
rect 107430 266782 107666 266868
rect 231814 266782 232050 267018
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 241382 266782 241618 267018
rect 244510 266782 244746 267018
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 61246 251142 61482 251378
rect 60878 249102 61114 249338
rect 59958 68902 60194 69138
rect 59590 68222 59826 68458
rect 61614 248422 61850 248658
rect 61062 72302 61298 72538
rect 62166 76532 62402 76618
rect 62166 76468 62252 76532
rect 62252 76468 62316 76532
rect 62316 76468 62402 76532
rect 62166 76382 62402 76468
rect 63638 68902 63874 69138
rect 64006 68222 64242 68458
rect 241198 266252 241434 266338
rect 241198 266188 241284 266252
rect 241284 266188 241348 266252
rect 241348 266188 241434 266252
rect 241198 266102 241434 266188
rect 201638 262702 201874 262938
rect 276894 44422 277130 44658
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 280022 266782 280258 267018
rect 279654 60742 279890 60978
rect 281310 77742 281546 77978
rect 281310 76532 281546 76618
rect 281310 76468 281396 76532
rect 281396 76468 281460 76532
rect 281460 76468 281546 76532
rect 281310 76382 281546 76468
rect 281310 72452 281546 72538
rect 281310 72388 281396 72452
rect 281396 72388 281460 72452
rect 281460 72388 281546 72452
rect 281310 72302 281546 72388
rect 281310 60892 281546 60978
rect 281310 60828 281396 60892
rect 281396 60828 281460 60892
rect 281460 60828 281546 60892
rect 281310 60742 281546 60828
rect 282046 248436 282282 248658
rect 282046 248422 282132 248436
rect 282132 248422 282196 248436
rect 282196 248422 282282 248436
rect 284254 262702 284490 262938
rect 282414 44422 282650 44658
rect 283334 251142 283570 251378
rect 283886 250462 284122 250698
rect 283334 72982 283570 73218
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 289590 267612 289826 267698
rect 289590 267548 289676 267612
rect 289676 267548 289740 267612
rect 289740 267548 289826 267612
rect 289590 267462 289826 267548
rect 291982 267612 292218 267698
rect 291982 267548 292068 267612
rect 292068 267548 292132 267612
rect 292132 267548 292218 267612
rect 291982 267462 292218 267548
rect 294558 266782 294794 267018
rect 299342 266932 299578 267018
rect 299342 266868 299428 266932
rect 299428 266868 299492 266932
rect 299492 266868 299578 266932
rect 299342 266782 299578 266868
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 320870 266932 321106 267018
rect 320870 266868 320956 266932
rect 320956 266868 321020 266932
rect 321020 266868 321106 266932
rect 320870 266782 321106 266868
rect 308910 266102 309146 266338
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 297870 77062 298106 77298
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288302 73132 288538 73218
rect 288302 73068 288388 73132
rect 288388 73068 288452 73132
rect 288452 73068 288538 73132
rect 288302 72982 288538 73068
rect 297870 73132 298106 73218
rect 297870 73068 297956 73132
rect 297956 73068 298020 73132
rect 298020 73068 298106 73132
rect 297870 72982 298106 73068
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 337982 266932 338218 267018
rect 337982 266868 338068 266932
rect 338068 266868 338132 266932
rect 338132 266868 338218 266932
rect 337982 266782 338218 266868
rect 328230 266102 328466 266338
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 318478 72302 318714 72538
rect 309094 71772 309330 71858
rect 309094 71708 309180 71772
rect 309180 71708 309244 71772
rect 309244 71708 309330 71772
rect 309094 71622 309330 71708
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 357302 266932 357538 267018
rect 357302 266868 357388 266932
rect 357388 266868 357452 266932
rect 357452 266868 357538 266932
rect 357302 266782 357538 266868
rect 347550 266102 347786 266338
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 337798 72302 338034 72538
rect 328414 71772 328650 71858
rect 328414 71708 328500 71772
rect 328500 71708 328564 71772
rect 328564 71708 328650 71772
rect 328414 71622 328650 71708
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 376806 266932 377042 267018
rect 376806 266868 376892 266932
rect 376892 266868 376956 266932
rect 376956 266868 377042 266932
rect 376806 266782 377042 266868
rect 366870 266102 367106 266338
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 357118 76382 357354 76618
rect 347734 75852 347970 75938
rect 347734 75788 347820 75852
rect 347820 75788 347884 75852
rect 347884 75788 347970 75852
rect 347734 75702 347970 75788
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 395942 266932 396178 267018
rect 395942 266868 396028 266932
rect 396028 266868 396092 266932
rect 396092 266868 396178 266932
rect 395942 266782 396178 266868
rect 386190 266102 386426 266338
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 376622 76532 376858 76618
rect 376622 76468 376708 76532
rect 376708 76468 376772 76532
rect 376772 76468 376858 76532
rect 376622 76382 376858 76468
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 357118 72302 357354 72538
rect 347734 71772 347970 71858
rect 347734 71708 347820 71772
rect 347820 71708 347884 71772
rect 347884 71708 347970 71772
rect 347734 71622 347970 71708
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 376438 72302 376674 72538
rect 378462 72452 378698 72538
rect 378462 72388 378548 72452
rect 378548 72388 378612 72452
rect 378612 72388 378698 72452
rect 378462 72302 378698 72388
rect 367054 71772 367290 71858
rect 367054 71708 367140 71772
rect 367140 71708 367204 71772
rect 367204 71708 367290 71772
rect 367054 71622 367290 71708
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 405510 266102 405746 266338
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 389686 76532 389922 76618
rect 389686 76468 389772 76532
rect 389772 76468 389836 76532
rect 389836 76468 389922 76532
rect 389686 76382 389922 76468
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 386190 72982 386426 73218
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 417470 266932 417706 267018
rect 417470 266868 417556 266932
rect 417556 266868 417620 266932
rect 417620 266868 417706 266932
rect 417470 266782 417706 266868
rect 424830 266102 425066 266338
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 405694 71622 405930 71858
rect 405694 69582 405930 69818
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 436790 266932 437026 267018
rect 436790 266868 436876 266932
rect 436876 266868 436940 266932
rect 436940 266868 437026 266932
rect 436790 266782 437026 266868
rect 444150 266102 444386 266338
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 415630 72452 415866 72538
rect 415630 72388 415716 72452
rect 415716 72388 415780 72452
rect 415780 72388 415866 72452
rect 415630 72302 415866 72388
rect 424830 71622 425066 71858
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 456110 266932 456346 267018
rect 456110 266868 456196 266932
rect 456196 266868 456260 266932
rect 456260 266868 456346 266932
rect 456110 266782 456346 266868
rect 463470 266102 463706 266338
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 437158 72452 437394 72538
rect 437158 72388 437244 72452
rect 437244 72388 437308 72452
rect 437308 72388 437394 72452
rect 437158 72302 437394 72388
rect 444150 72452 444386 72538
rect 444150 72388 444236 72452
rect 444236 72388 444300 72452
rect 444300 72388 444386 72452
rect 444150 72302 444386 72388
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 475430 266932 475666 267018
rect 475430 266868 475516 266932
rect 475516 266868 475580 266932
rect 475580 266868 475666 266932
rect 475430 266782 475666 266868
rect 482790 266102 483026 266338
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 453902 71772 454138 71858
rect 453902 71708 453988 71772
rect 453988 71708 454052 71772
rect 454052 71708 454138 71772
rect 453902 71622 454138 71708
rect 463470 71772 463706 71858
rect 463470 71708 463556 71772
rect 463556 71708 463620 71772
rect 463620 71708 463706 71772
rect 463470 71622 463706 71708
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 492726 266932 492962 267018
rect 492726 266868 492812 266932
rect 492812 266868 492876 266932
rect 492876 266868 492962 266932
rect 492726 266782 492962 266868
rect 502110 266102 502346 266338
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 475246 72452 475482 72538
rect 475246 72388 475332 72452
rect 475332 72388 475396 72452
rect 475396 72388 475482 72452
rect 475246 72302 475482 72388
rect 476166 72452 476402 72538
rect 476166 72388 476252 72452
rect 476252 72388 476316 72452
rect 476316 72388 476402 72452
rect 476166 72302 476402 72388
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 511862 266932 512098 267018
rect 511862 266868 511948 266932
rect 511948 266868 512012 266932
rect 512012 266868 512098 266932
rect 511862 266782 512098 266868
rect 521430 266102 521666 266338
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 494750 77212 494986 77298
rect 494750 77148 494836 77212
rect 494836 77148 494900 77212
rect 494900 77148 494986 77212
rect 494750 77062 494986 77148
rect 500638 76382 500874 76618
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 502294 71772 502530 71858
rect 502294 71708 502380 71772
rect 502380 71708 502444 71772
rect 502444 71708 502530 71772
rect 502294 71622 502530 71708
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 533758 267462 533994 267698
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 511678 71772 511914 71858
rect 511678 71708 511764 71772
rect 511764 71708 511828 71772
rect 511828 71708 511914 71772
rect 511678 71622 511914 71708
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 552526 73132 552762 73218
rect 552526 73068 552612 73132
rect 552612 73068 552676 73132
rect 552676 73068 552762 73132
rect 552526 72982 552762 73068
rect 553446 73132 553682 73218
rect 553446 73068 553532 73132
rect 553532 73068 553596 73132
rect 553596 73068 553682 73132
rect 553446 72982 553682 73068
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 580678 76382 580914 76618
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 580310 72982 580546 73218
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect 109044 267420 118932 267740
rect 109044 267060 109364 267420
rect 107388 267018 109364 267060
rect 107388 266782 107430 267018
rect 107666 266782 109364 267018
rect 107388 266740 109364 266782
rect 118612 267060 118932 267420
rect 132412 267420 142484 267740
rect 132412 267060 132732 267420
rect 118612 266740 132732 267060
rect 142164 267060 142484 267420
rect 151732 267420 161804 267740
rect 151732 267060 152052 267420
rect 142164 266740 152052 267060
rect 161484 267060 161804 267420
rect 171052 267420 181124 267740
rect 171052 267060 171372 267420
rect 161484 266740 171372 267060
rect 180804 267060 181124 267420
rect 190372 267420 200260 267740
rect 190372 267060 190692 267420
rect 180804 266740 190692 267060
rect 199940 267060 200260 267420
rect 205644 267420 225284 267740
rect 205644 267060 205964 267420
rect 199940 266740 205964 267060
rect 224964 267060 225284 267420
rect 253852 267420 260980 267740
rect 289548 267698 292260 267740
rect 289548 267462 289590 267698
rect 289826 267462 291982 267698
rect 292218 267462 292260 267698
rect 289548 267420 292260 267462
rect 524332 267698 534036 267740
rect 524332 267462 533758 267698
rect 533994 267462 534036 267698
rect 524332 267420 534036 267462
rect 253852 267060 254172 267420
rect 224964 267018 232092 267060
rect 224964 266782 231814 267018
rect 232050 266782 232092 267018
rect 224964 266740 232092 266782
rect 241340 267018 241660 267060
rect 241340 266782 241382 267018
rect 241618 266782 241660 267018
rect 241340 266380 241660 266782
rect 244468 267018 254172 267060
rect 244468 266782 244510 267018
rect 244746 266782 254172 267018
rect 244468 266740 254172 266782
rect 260660 267060 260980 267420
rect 260660 267018 280300 267060
rect 260660 266782 280022 267018
rect 280258 266782 280300 267018
rect 260660 266740 280300 266782
rect 294516 267018 299620 267060
rect 294516 266782 294558 267018
rect 294794 266782 299342 267018
rect 299578 266782 299620 267018
rect 294516 266740 299620 266782
rect 311812 267018 321148 267060
rect 311812 266782 320870 267018
rect 321106 266782 321148 267018
rect 311812 266740 321148 266782
rect 331132 267018 338260 267060
rect 331132 266782 337982 267018
rect 338218 266782 338260 267018
rect 331132 266740 338260 266782
rect 350452 267018 357580 267060
rect 350452 266782 357302 267018
rect 357538 266782 357580 267018
rect 350452 266740 357580 266782
rect 369772 267018 377084 267060
rect 369772 266782 376806 267018
rect 377042 266782 377084 267018
rect 369772 266740 377084 266782
rect 389092 267018 396220 267060
rect 389092 266782 395942 267018
rect 396178 266782 396220 267018
rect 389092 266740 396220 266782
rect 408412 267018 417748 267060
rect 408412 266782 417470 267018
rect 417706 266782 417748 267018
rect 408412 266740 417748 266782
rect 427732 267018 437068 267060
rect 427732 266782 436790 267018
rect 437026 266782 437068 267018
rect 427732 266740 437068 266782
rect 447052 267018 456388 267060
rect 447052 266782 456110 267018
rect 456346 266782 456388 267018
rect 447052 266740 456388 266782
rect 466372 267018 475708 267060
rect 466372 266782 475430 267018
rect 475666 266782 475708 267018
rect 466372 266740 475708 266782
rect 485692 267018 493004 267060
rect 485692 266782 492726 267018
rect 492962 266782 493004 267018
rect 485692 266740 493004 266782
rect 505012 267018 512140 267060
rect 505012 266782 511862 267018
rect 512098 266782 512140 267018
rect 505012 266740 512140 266782
rect 311812 266380 312132 266740
rect 331132 266380 331452 266740
rect 350452 266380 350772 266740
rect 369772 266380 370092 266740
rect 389092 266380 389412 266740
rect 408412 266380 408732 266740
rect 427732 266380 428052 266740
rect 447052 266380 447372 266740
rect 466372 266380 466692 266740
rect 485692 266380 486012 266740
rect 505012 266380 505332 266740
rect 524332 266380 524652 267420
rect 241156 266338 241660 266380
rect 241156 266102 241198 266338
rect 241434 266102 241660 266338
rect 241156 266060 241660 266102
rect 308868 266338 312132 266380
rect 308868 266102 308910 266338
rect 309146 266102 312132 266338
rect 308868 266060 312132 266102
rect 328188 266338 331452 266380
rect 328188 266102 328230 266338
rect 328466 266102 331452 266338
rect 328188 266060 331452 266102
rect 347508 266338 350772 266380
rect 347508 266102 347550 266338
rect 347786 266102 350772 266338
rect 347508 266060 350772 266102
rect 366828 266338 370092 266380
rect 366828 266102 366870 266338
rect 367106 266102 370092 266338
rect 366828 266060 370092 266102
rect 386148 266338 389412 266380
rect 386148 266102 386190 266338
rect 386426 266102 389412 266338
rect 386148 266060 389412 266102
rect 405468 266338 408732 266380
rect 405468 266102 405510 266338
rect 405746 266102 408732 266338
rect 405468 266060 408732 266102
rect 424788 266338 428052 266380
rect 424788 266102 424830 266338
rect 425066 266102 428052 266338
rect 424788 266060 428052 266102
rect 444108 266338 447372 266380
rect 444108 266102 444150 266338
rect 444386 266102 447372 266338
rect 444108 266060 447372 266102
rect 463428 266338 466692 266380
rect 463428 266102 463470 266338
rect 463706 266102 466692 266338
rect 463428 266060 466692 266102
rect 482748 266338 486012 266380
rect 482748 266102 482790 266338
rect 483026 266102 486012 266338
rect 482748 266060 486012 266102
rect 502068 266338 505332 266380
rect 502068 266102 502110 266338
rect 502346 266102 505332 266338
rect 502068 266060 505332 266102
rect 521388 266338 524652 266380
rect 521388 266102 521430 266338
rect 521666 266102 524652 266338
rect 521388 266060 524652 266102
rect 201596 262938 284532 262980
rect 201596 262702 201638 262938
rect 201874 262702 284254 262938
rect 284490 262702 284532 262938
rect 201596 262660 284532 262702
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect 74636 253140 83236 253460
rect 74636 251420 74956 253140
rect 82916 252100 83236 253140
rect 92300 253140 100532 253460
rect 92300 252780 92620 253140
rect 91196 252460 92620 252780
rect 100212 252780 100532 253140
rect 110332 253140 112676 253460
rect 110332 252780 110652 253140
rect 100212 252460 102188 252780
rect 82916 251780 85076 252100
rect 84756 251420 85076 251780
rect 91196 251420 91516 252460
rect 101868 252100 102188 252460
rect 110148 252460 110652 252780
rect 110148 252100 110468 252460
rect 101868 251780 110468 252100
rect 112356 252100 112676 253140
rect 121556 253140 130892 253460
rect 112356 251780 120956 252100
rect 61204 251378 74956 251420
rect 61204 251142 61246 251378
rect 61482 251142 74956 251378
rect 61204 251100 74956 251142
rect 77028 251100 84340 251420
rect 84756 251100 91516 251420
rect 99844 251100 100900 251420
rect 101868 251100 102372 251780
rect 120636 251420 120956 251780
rect 121556 251420 121876 253140
rect 104076 251100 111204 251420
rect 120636 251100 121876 251420
rect 130572 251420 130892 253140
rect 142164 253140 155364 253460
rect 131676 251780 140276 252100
rect 131676 251420 131996 251780
rect 130572 251100 131996 251420
rect 139956 251420 140276 251780
rect 142164 251420 142484 253140
rect 155044 252100 155364 253140
rect 161484 253140 174684 253460
rect 155044 251780 159780 252100
rect 159460 251420 159780 251780
rect 161484 251420 161804 253140
rect 174364 252100 174684 253140
rect 189084 253140 198604 253460
rect 174364 251780 179100 252100
rect 178780 251420 179100 251780
rect 189084 251420 189404 253140
rect 139956 251100 142484 251420
rect 150444 251100 159044 251420
rect 159460 251100 161804 251420
rect 169764 251100 178364 251420
rect 178780 251100 184436 251420
rect 67460 249740 74772 250060
rect 67460 249380 67780 249740
rect 60836 249338 67780 249380
rect 60836 249102 60878 249338
rect 61114 249102 67780 249338
rect 60836 249060 67780 249102
rect 74452 249380 74772 249740
rect 77028 249380 77348 251100
rect 81076 250420 82500 250740
rect 74452 249060 77348 249380
rect 77764 249740 79188 250060
rect 77764 248700 78084 249740
rect 78868 249380 79188 249740
rect 81076 249380 81396 250420
rect 78868 249060 81396 249380
rect 82180 249380 82500 250420
rect 84020 250060 84340 251100
rect 99844 250740 100164 251100
rect 90644 250420 92436 250740
rect 90644 250060 90964 250420
rect 84020 249740 90964 250060
rect 92116 250060 92436 250420
rect 93588 250420 100164 250740
rect 100580 250740 100900 251100
rect 104076 250740 104396 251100
rect 100580 250420 104396 250740
rect 110884 250740 111204 251100
rect 110884 250420 111756 250740
rect 93588 250060 93908 250420
rect 111436 250060 111756 250420
rect 121004 250420 129052 250740
rect 121004 250060 121324 250420
rect 92116 249740 93908 250060
rect 100212 249740 101268 250060
rect 82180 249060 84156 249380
rect 61572 248658 78084 248700
rect 61572 248422 61614 248658
rect 61850 248422 78084 248658
rect 61572 248380 78084 248422
rect 83836 248700 84156 249060
rect 100212 248700 100532 249740
rect 100948 249380 101268 249740
rect 102420 249740 103660 250060
rect 102420 249380 102740 249740
rect 100948 249060 102740 249380
rect 83836 248380 100532 248700
rect 103340 248700 103660 249740
rect 106836 249740 110836 250060
rect 111436 249740 112308 250060
rect 106836 248700 107156 249740
rect 103340 248380 107156 248700
rect 110516 248700 110836 249740
rect 111988 249380 112308 249740
rect 116956 249740 121324 250060
rect 128732 250060 129052 250420
rect 140324 250420 148004 250740
rect 140324 250060 140644 250420
rect 128732 249740 131628 250060
rect 116956 249380 117276 249740
rect 131308 249380 131628 249740
rect 136276 249740 140644 250060
rect 136276 249380 136596 249740
rect 147684 249380 148004 250420
rect 150444 249380 150764 251100
rect 158724 250740 159044 251100
rect 158724 250420 167324 250740
rect 167004 249380 167324 250420
rect 169764 249380 170084 251100
rect 178044 250740 178364 251100
rect 184116 250740 184436 251100
rect 188532 251100 189404 251420
rect 198284 251420 198604 253140
rect 209876 253140 219212 253460
rect 209876 251420 210196 253140
rect 218892 251420 219212 253140
rect 229196 253140 238532 253460
rect 229196 251420 229516 253140
rect 238212 251420 238532 253140
rect 248516 253140 257852 253460
rect 248516 251420 248836 253140
rect 257532 251420 257852 253140
rect 198284 251100 210196 251420
rect 210612 251100 215532 251420
rect 218892 251100 229516 251420
rect 229932 251100 234852 251420
rect 238212 251100 248836 251420
rect 249252 251100 254172 251420
rect 257532 251378 283612 251420
rect 257532 251142 283334 251378
rect 283570 251142 283612 251378
rect 257532 251100 283612 251142
rect 188532 250740 188852 251100
rect 178044 250420 179836 250740
rect 184116 250420 188852 250740
rect 189268 250420 196948 250740
rect 179516 250060 179836 250420
rect 189268 250060 189588 250420
rect 179516 249740 189588 250060
rect 196628 249380 196948 250420
rect 209508 250060 210012 250740
rect 210612 250060 210932 251100
rect 209508 249740 210932 250060
rect 215212 250060 215532 251100
rect 222204 250420 229332 250740
rect 222204 250060 222524 250420
rect 215212 249740 219396 250060
rect 209508 249380 209828 249740
rect 111988 249060 117276 249380
rect 121188 249060 124820 249380
rect 131308 249060 136596 249380
rect 140508 249060 144324 249380
rect 147684 249060 150764 249380
rect 159828 249060 163644 249380
rect 167004 249060 170084 249380
rect 179148 249060 182780 249380
rect 196628 249060 209828 249380
rect 219076 249380 219396 249740
rect 222020 249740 222524 250060
rect 229012 250060 229332 250420
rect 229932 250060 230252 251100
rect 229012 249740 230252 250060
rect 234532 250060 234852 251100
rect 241524 250420 248652 250740
rect 241524 250060 241844 250420
rect 234532 249740 238716 250060
rect 222020 249380 222340 249740
rect 219076 249060 222340 249380
rect 238396 249380 238716 249740
rect 241340 249740 241844 250060
rect 248332 250060 248652 250420
rect 249252 250060 249572 251100
rect 248332 249740 249572 250060
rect 253852 250060 254172 251100
rect 273172 250698 284164 250740
rect 273172 250462 283886 250698
rect 284122 250462 284164 250698
rect 273172 250420 284164 250462
rect 273172 250060 273492 250420
rect 253852 249740 258036 250060
rect 241340 249380 241660 249740
rect 238396 249060 241660 249380
rect 257716 249380 258036 249740
rect 262868 249740 273492 250060
rect 262868 249380 263188 249740
rect 257716 249060 263188 249380
rect 121188 248700 121508 249060
rect 110516 248380 121508 248700
rect 124500 248700 124820 249060
rect 140508 248700 140828 249060
rect 124500 248380 140828 248700
rect 144004 248700 144324 249060
rect 159828 248700 160148 249060
rect 144004 248380 160148 248700
rect 163324 248700 163644 249060
rect 179148 248700 179468 249060
rect 163324 248380 179468 248700
rect 182460 248700 182780 249060
rect 182460 248658 282324 248700
rect 182460 248422 282046 248658
rect 282282 248422 282324 248658
rect 182460 248380 282324 248422
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect 3244 79338 9820 79380
rect 3244 79102 3286 79338
rect 3522 79102 9820 79338
rect 3244 79060 9820 79102
rect 9500 78700 9820 79060
rect 12260 79060 19388 79380
rect 22564 79338 29140 79380
rect 22564 79102 22606 79338
rect 22842 79102 28862 79338
rect 29098 79102 29140 79338
rect 22564 79060 29140 79102
rect 41884 79338 47172 79380
rect 41884 79102 41926 79338
rect 42162 79102 47172 79338
rect 41884 79060 47172 79102
rect 12260 78700 12580 79060
rect 9500 78380 12580 78700
rect 19068 78700 19388 79060
rect 46852 78700 47172 79060
rect 50900 79060 60190 79380
rect 50900 78700 51220 79060
rect 19068 78380 19756 78700
rect 46852 78380 51220 78700
rect 59870 78700 60190 79060
rect 59870 78380 70724 78700
rect 19436 77978 19756 78380
rect 19436 77742 19478 77978
rect 19714 77742 19756 77978
rect 19436 77700 19756 77742
rect 70404 78020 70724 78380
rect 88620 78380 90780 78700
rect 88620 78020 88940 78380
rect 90460 78020 90780 78380
rect 95060 78380 104948 78700
rect 95060 78020 95380 78380
rect 70404 77700 88940 78020
rect 89356 77340 89860 78020
rect 90460 77700 95380 78020
rect 104628 78020 104948 78380
rect 107940 78380 110100 78700
rect 107940 78020 108260 78380
rect 109780 78020 110100 78380
rect 114380 78380 124268 78700
rect 114380 78020 114700 78380
rect 104628 77700 108260 78020
rect 108676 77340 109180 78020
rect 109780 77700 114700 78020
rect 123948 78020 124268 78380
rect 127260 78380 129420 78700
rect 127260 78020 127580 78380
rect 129100 78020 129420 78380
rect 133700 78380 143588 78700
rect 133700 78020 134020 78380
rect 123948 77700 127580 78020
rect 127996 77340 128500 78020
rect 129100 77700 134020 78020
rect 143268 78020 143588 78380
rect 146580 78380 148740 78700
rect 146580 78020 146900 78380
rect 148420 78020 148740 78380
rect 153020 78380 162908 78700
rect 153020 78020 153340 78380
rect 143268 77700 146900 78020
rect 147316 77340 147820 78020
rect 148420 77700 153340 78020
rect 162588 78020 162908 78380
rect 165900 78380 168060 78700
rect 165900 78020 166220 78380
rect 167740 78020 168060 78380
rect 172340 78380 182228 78700
rect 172340 78020 172660 78380
rect 162588 77700 166220 78020
rect 166636 77340 167140 78020
rect 167740 77700 172660 78020
rect 181908 78020 182228 78380
rect 185220 78380 187380 78700
rect 185220 78020 185540 78380
rect 187060 78020 187380 78380
rect 191660 78380 201548 78700
rect 191660 78020 191980 78380
rect 181908 77700 185540 78020
rect 185956 77340 186460 78020
rect 187060 77700 191980 78020
rect 201228 78020 201548 78380
rect 204540 78380 206700 78700
rect 204540 78020 204860 78380
rect 206380 78020 206700 78380
rect 210980 78380 220868 78700
rect 210980 78020 211300 78380
rect 201228 77700 204860 78020
rect 205276 77340 205780 78020
rect 206380 77700 211300 78020
rect 220548 78020 220868 78380
rect 223860 78380 226020 78700
rect 223860 78020 224180 78380
rect 225700 78020 226020 78380
rect 230300 78380 240188 78700
rect 230300 78020 230620 78380
rect 220548 77700 224180 78020
rect 224596 77340 225100 78020
rect 225700 77700 230620 78020
rect 239868 78020 240188 78380
rect 243180 78380 245340 78700
rect 243180 78020 243500 78380
rect 245020 78020 245340 78380
rect 249620 78380 259508 78700
rect 249620 78020 249940 78380
rect 239868 77700 243500 78020
rect 243916 77340 244420 78020
rect 245020 77700 249940 78020
rect 259188 78020 259508 78380
rect 262500 78380 264660 78700
rect 262500 78020 262820 78380
rect 259188 77700 262820 78020
rect 264340 78020 264660 78380
rect 272252 78380 281588 78700
rect 272252 78020 272572 78380
rect 264340 77700 272572 78020
rect 74452 77020 89860 77340
rect 62124 76618 67780 76660
rect 62124 76382 62166 76618
rect 62402 76382 67780 76618
rect 62124 76340 67780 76382
rect 67460 75980 67780 76340
rect 74452 75980 74772 77020
rect 89540 76660 89860 77020
rect 95244 77020 109180 77340
rect 95244 76660 95564 77020
rect 89540 76340 95564 76660
rect 108860 76660 109180 77020
rect 114564 77020 128500 77340
rect 114564 76660 114884 77020
rect 108860 76340 114884 76660
rect 128180 76660 128500 77020
rect 133884 77020 147820 77340
rect 133884 76660 134204 77020
rect 128180 76340 134204 76660
rect 147500 76660 147820 77020
rect 153204 77020 167140 77340
rect 153204 76660 153524 77020
rect 147500 76340 153524 76660
rect 166820 76660 167140 77020
rect 172524 77020 186460 77340
rect 172524 76660 172844 77020
rect 166820 76340 172844 76660
rect 186140 76660 186460 77020
rect 191844 77020 205780 77340
rect 191844 76660 192164 77020
rect 186140 76340 192164 76660
rect 205460 76660 205780 77020
rect 211164 77020 225100 77340
rect 211164 76660 211484 77020
rect 205460 76340 211484 76660
rect 224780 76660 225100 77020
rect 230484 77020 244420 77340
rect 230484 76660 230804 77020
rect 224780 76340 230804 76660
rect 244100 76660 244420 77020
rect 249804 77020 263372 77340
rect 249804 76660 250124 77020
rect 244100 76340 250124 76660
rect 67460 75660 74772 75980
rect 263052 75300 263372 77020
rect 272988 76660 273492 78020
rect 281268 77978 281588 78380
rect 281268 77742 281310 77978
rect 281546 77742 281588 77978
rect 281268 77700 281588 77742
rect 398476 77700 409284 78020
rect 297828 77298 299620 77340
rect 297828 77062 297870 77298
rect 298106 77062 299620 77298
rect 297828 77020 299620 77062
rect 299300 76660 299620 77020
rect 337756 77020 341020 77340
rect 270228 76618 281588 76660
rect 270228 76382 281310 76618
rect 281546 76382 281588 76618
rect 270228 76340 281588 76382
rect 299300 76340 309188 76660
rect 270228 75300 270548 76340
rect 308868 75980 309188 76340
rect 318436 76340 321516 76660
rect 318436 75980 318756 76340
rect 308868 75660 318756 75980
rect 321196 75980 321516 76340
rect 337756 75980 338076 77020
rect 321196 75660 338076 75980
rect 340700 75980 341020 77020
rect 398476 76660 398796 77700
rect 408964 77340 409284 77700
rect 417244 77700 418300 78020
rect 417244 77340 417564 77700
rect 408964 77020 417564 77340
rect 357076 76618 360156 76660
rect 357076 76382 357118 76618
rect 357354 76382 360156 76618
rect 357076 76340 360156 76382
rect 359836 75980 360156 76340
rect 376396 76618 377056 76660
rect 376396 76382 376622 76618
rect 376858 76382 377056 76618
rect 376396 76340 377056 76382
rect 389644 76618 398796 76660
rect 389644 76382 389686 76618
rect 389922 76382 398796 76618
rect 389644 76340 398796 76382
rect 417980 76660 418300 77700
rect 427548 77340 428052 78020
rect 437116 77340 437620 78020
rect 427548 77020 437620 77340
rect 427548 76660 427868 77020
rect 417980 76340 427868 76660
rect 437300 76660 437620 77020
rect 446868 76660 447372 78020
rect 456436 77700 476260 78020
rect 456436 76660 456756 77700
rect 437300 76340 456756 76660
rect 475940 76660 476260 77700
rect 485508 77340 486012 78020
rect 504828 77700 505884 78020
rect 485508 77298 495028 77340
rect 485508 77062 494750 77298
rect 494986 77062 495028 77298
rect 485508 77020 495028 77062
rect 485508 76660 485828 77020
rect 504828 76660 505148 77700
rect 505564 77340 505884 77700
rect 513844 77700 514900 78020
rect 513844 77340 514164 77700
rect 505564 77020 514164 77340
rect 475940 76340 485828 76660
rect 500596 76618 505148 76660
rect 500596 76382 500638 76618
rect 500874 76382 505148 76618
rect 500596 76340 505148 76382
rect 514580 76660 514900 77700
rect 524148 77700 534772 78020
rect 524148 76660 524468 77700
rect 534452 77340 534772 77700
rect 552484 77700 553540 78020
rect 552484 77340 552804 77700
rect 534452 77020 552804 77340
rect 514580 76340 524468 76660
rect 553220 76660 553540 77700
rect 562788 77700 567340 78020
rect 562788 76660 563108 77700
rect 553220 76340 563108 76660
rect 567020 76660 567340 77700
rect 567020 76618 580956 76660
rect 567020 76382 580678 76618
rect 580914 76382 580956 76618
rect 567020 76340 580956 76382
rect 376396 75980 376716 76340
rect 340700 75938 348012 75980
rect 340700 75702 347734 75938
rect 347970 75702 348012 75938
rect 340700 75660 348012 75702
rect 359836 75660 376716 75980
rect 263052 74980 270548 75300
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect 69852 72940 87284 73260
rect 69852 72580 70172 72940
rect 61020 72538 70172 72580
rect 61020 72302 61062 72538
rect 61298 72302 70172 72538
rect 61020 72260 70172 72302
rect 79788 71580 80292 72940
rect 86964 71900 87284 72940
rect 99476 72940 106604 73260
rect 99476 71900 99796 72940
rect 86964 71580 87468 71900
rect 87148 69180 87468 71580
rect 96164 71580 99796 71900
rect 106284 71900 106604 72940
rect 118796 72940 125924 73260
rect 118796 71900 119116 72940
rect 106284 71580 106788 71900
rect 96164 69180 96484 71580
rect 59916 69138 63916 69180
rect 59916 68902 59958 69138
rect 60194 68902 63638 69138
rect 63874 68902 63916 69138
rect 59916 68860 63916 68902
rect 87148 68860 96484 69180
rect 106468 69180 106788 71580
rect 115484 71580 119116 71900
rect 125604 71900 125924 72940
rect 138116 72940 145244 73260
rect 138116 71900 138436 72940
rect 125604 71580 126108 71900
rect 115484 69180 115804 71580
rect 106468 68860 115804 69180
rect 125788 69180 126108 71580
rect 134804 71580 138436 71900
rect 144924 71900 145244 72940
rect 157436 72940 164564 73260
rect 157436 71900 157756 72940
rect 144924 71580 145428 71900
rect 134804 69180 135124 71580
rect 125788 68860 135124 69180
rect 145108 69180 145428 71580
rect 154124 71580 157756 71900
rect 164244 71900 164564 72940
rect 176756 72940 183884 73260
rect 176756 71900 177076 72940
rect 164244 71580 164748 71900
rect 154124 69180 154444 71580
rect 145108 68860 154444 69180
rect 164428 69180 164748 71580
rect 173444 71580 177076 71900
rect 183564 71900 183884 72940
rect 196076 72940 203204 73260
rect 196076 71900 196396 72940
rect 183564 71580 184068 71900
rect 173444 69180 173764 71580
rect 164428 68860 173764 69180
rect 183748 69180 184068 71580
rect 192764 71580 196396 71900
rect 202884 71900 203204 72940
rect 215396 72940 222524 73260
rect 215396 71900 215716 72940
rect 202884 71580 203388 71900
rect 192764 69180 193084 71580
rect 183748 68860 193084 69180
rect 203068 69180 203388 71580
rect 212084 71580 215716 71900
rect 222204 71900 222524 72940
rect 234716 72940 241844 73260
rect 234716 71900 235036 72940
rect 222204 71580 222708 71900
rect 212084 69180 212404 71580
rect 203068 68860 212404 69180
rect 222388 69180 222708 71580
rect 231404 71580 235036 71900
rect 241524 71900 241844 72940
rect 254036 72940 265764 73260
rect 283292 73218 288580 73260
rect 283292 72982 283334 73218
rect 283570 72982 288302 73218
rect 288538 72982 288580 73218
rect 283292 72940 288580 72982
rect 297828 73218 299620 73260
rect 297828 72982 297870 73218
rect 298106 72982 299620 73218
rect 297828 72940 299620 72982
rect 386148 73218 389228 73260
rect 386148 72982 386190 73218
rect 386426 72982 389228 73218
rect 386148 72940 389228 72982
rect 254036 71900 254356 72940
rect 241524 71580 242028 71900
rect 231404 69180 231724 71580
rect 222388 68860 231724 69180
rect 241708 69180 242028 71580
rect 250724 71580 254356 71900
rect 265444 71900 265764 72940
rect 299300 72580 299620 72940
rect 273172 72538 281588 72580
rect 273172 72302 281310 72538
rect 281546 72302 281588 72538
rect 273172 72260 281588 72302
rect 299300 72260 309188 72580
rect 318436 72538 321516 72580
rect 318436 72302 318478 72538
rect 318714 72302 321516 72538
rect 318436 72260 321516 72302
rect 337756 72538 340836 72580
rect 337756 72302 337798 72538
rect 338034 72302 340836 72538
rect 337756 72260 340836 72302
rect 357076 72538 360156 72580
rect 357076 72302 357118 72538
rect 357354 72302 360156 72538
rect 357076 72260 360156 72302
rect 376396 72538 378740 72580
rect 376396 72302 376438 72538
rect 376674 72302 378462 72538
rect 378698 72302 378740 72538
rect 376396 72260 378740 72302
rect 273172 71900 273492 72260
rect 265444 71580 273492 71900
rect 308868 71900 309188 72260
rect 321196 71900 321516 72260
rect 340516 71900 340836 72260
rect 359836 71900 360156 72260
rect 388908 71900 389228 72940
rect 514396 72940 528700 73260
rect 389644 72260 398428 72580
rect 389644 71900 389964 72260
rect 308868 71858 309372 71900
rect 308868 71622 309094 71858
rect 309330 71622 309372 71858
rect 308868 71580 309372 71622
rect 321196 71858 328692 71900
rect 321196 71622 328414 71858
rect 328650 71622 328692 71858
rect 321196 71580 328692 71622
rect 340516 71858 348012 71900
rect 340516 71622 347734 71858
rect 347970 71622 348012 71858
rect 340516 71580 348012 71622
rect 359836 71858 367332 71900
rect 359836 71622 367054 71858
rect 367290 71622 367332 71858
rect 359836 71580 367332 71622
rect 388908 71580 389964 71900
rect 398108 71900 398428 72260
rect 414852 72538 415908 72580
rect 414852 72302 415630 72538
rect 415866 72302 415908 72538
rect 414852 72260 415908 72302
rect 424972 72538 437436 72580
rect 424972 72302 437158 72538
rect 437394 72302 437436 72538
rect 424972 72260 437436 72302
rect 444108 72538 444796 72580
rect 444108 72302 444150 72538
rect 444386 72302 444796 72538
rect 444108 72260 444796 72302
rect 398108 71858 405972 71900
rect 398108 71622 405694 71858
rect 405930 71622 405972 71858
rect 398108 71580 405972 71622
rect 250724 69180 251044 71580
rect 414852 69860 415172 72260
rect 424972 71900 425292 72260
rect 424632 71858 425292 71900
rect 424632 71622 424830 71858
rect 425066 71622 425292 71858
rect 424632 71580 425292 71622
rect 444476 71900 444796 72260
rect 472996 72538 475524 72580
rect 472996 72302 475246 72538
rect 475482 72302 475524 72538
rect 472996 72260 475524 72302
rect 476124 72538 485276 72580
rect 476124 72302 476166 72538
rect 476402 72302 485276 72538
rect 476124 72260 485276 72302
rect 472996 71900 473316 72260
rect 444476 71858 454180 71900
rect 444476 71622 453902 71858
rect 454138 71622 454180 71858
rect 444476 71580 454180 71622
rect 463428 71858 473316 71900
rect 463428 71622 463470 71858
rect 463706 71622 473316 71858
rect 463428 71580 473316 71622
rect 484956 71900 485276 72260
rect 486244 72260 495028 72580
rect 486244 71900 486564 72260
rect 484956 71580 486564 71900
rect 494708 71900 495028 72260
rect 514396 71900 514716 72940
rect 494708 71858 502572 71900
rect 494708 71622 502294 71858
rect 502530 71622 502572 71858
rect 494708 71580 502572 71622
rect 511636 71858 514716 71900
rect 511636 71622 511678 71858
rect 511914 71622 514716 71858
rect 511636 71580 514716 71622
rect 528380 71900 528700 72940
rect 534452 73218 552804 73260
rect 534452 72982 552526 73218
rect 552762 72982 552804 73218
rect 534452 72940 552804 72982
rect 553404 73218 563108 73260
rect 553404 72982 553446 73218
rect 553682 72982 563108 73218
rect 553404 72940 563108 72982
rect 534452 71900 534772 72940
rect 528380 71580 534772 71900
rect 562788 71900 563108 72940
rect 566836 73218 580588 73260
rect 566836 72982 580310 73218
rect 580546 72982 580588 73218
rect 566836 72940 580588 72982
rect 566836 71900 567156 72940
rect 562788 71580 567156 71900
rect 405652 69818 415172 69860
rect 405652 69582 405694 69818
rect 405930 69582 415172 69818
rect 405652 69540 415172 69582
rect 241708 68860 251044 69180
rect 59548 68458 64284 68500
rect 59548 68222 59590 68458
rect 59826 68222 64006 68458
rect 64242 68222 64284 68458
rect 59548 68180 64284 68222
rect 279612 60978 281588 61020
rect 279612 60742 279654 60978
rect 279890 60742 281310 60978
rect 281546 60742 281588 60978
rect 279612 60700 281588 60742
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect 276852 44658 282692 44700
rect 276852 44422 276894 44658
rect 277130 44422 282414 44658
rect 282650 44422 282692 44658
rect 276852 44380 282692 44422
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 591900 -7506 592500 -7504
use tinyriscv  mprj
timestamp 1609751852
transform 1 0 62000 0 1 43200
box 0 0 219661 221805
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew signal input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew signal input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew signal input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew signal input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew signal input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew signal input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew signal input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew signal input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew signal input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew signal input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew signal input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew signal input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew signal input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew signal input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew signal input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew signal input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew signal input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew signal input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew signal input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew signal input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew signal input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew signal input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew signal input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew signal input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew signal input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew signal input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew signal input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew signal input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew signal input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew signal tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew signal tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew signal tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew signal tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew signal tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew signal tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew signal tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew signal tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew signal tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew signal tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew signal tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew signal tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew signal tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew signal tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew signal tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew signal tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew signal tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew signal tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew signal tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew signal tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew signal tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew signal tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew signal tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew signal tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew signal tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew signal tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew signal tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew signal tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew signal tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew signal tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew signal tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew signal tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew signal tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew signal tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew signal tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew signal tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew signal tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew signal tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew signal tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew signal tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew signal tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew signal tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew signal tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew signal tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew signal tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew signal tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew signal tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew signal tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew signal tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew signal tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew signal tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew signal tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew signal tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew signal tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew signal tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew signal tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew signal tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew signal tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew signal tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew signal tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew signal tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew signal tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew signal tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew signal tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew signal tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew signal tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew signal tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew signal tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew signal tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew signal tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew signal tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew signal tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew signal tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew signal tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew signal tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew signal tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew signal tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew signal tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew signal tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew signal tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew signal tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew signal tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew signal tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew signal tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew signal tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew signal tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew signal tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew signal tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew signal tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew signal tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew signal tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew signal tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew signal tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew signal tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew signal tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew signal tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew signal tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew signal tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew signal tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew signal tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew signal tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew signal tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew signal tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew signal tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew signal tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew signal tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew signal tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew signal tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew signal tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew signal tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew signal tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew signal tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew signal tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew signal tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew signal tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew signal tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew signal tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew signal tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew signal tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew signal tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew signal tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew signal tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew signal tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew signal tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew signal tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew signal tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew signal tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew signal tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew signal tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew signal tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew signal tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew signal tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew signal tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew signal tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew signal tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew signal tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew signal tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew signal tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew signal tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew signal tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew signal tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew signal tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew signal tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew signal tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew signal tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew signal tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew signal tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew signal tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew signal tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew signal tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew signal tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew signal tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew signal tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew signal tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew signal tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew signal tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew signal tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew signal tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew signal tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew signal tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew signal tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew signal tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew signal tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew signal tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew signal tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew signal tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew signal tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew signal tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew signal tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew signal tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew signal tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew signal tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew signal tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew signal tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew signal tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew signal tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew signal tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew signal tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew signal tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew signal tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew signal tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew signal tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew signal tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew signal tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew signal tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew signal input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew signal input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew signal input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew signal input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew signal input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew signal input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew signal input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew signal input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew signal input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew signal input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew signal input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew signal input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew signal input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew signal input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew signal input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew signal input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew signal input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew signal input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew signal input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew signal input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew signal input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew signal input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew signal input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew signal input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew signal input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew signal input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew signal input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew signal input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew signal input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew signal input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew signal input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew signal input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew signal input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew signal input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew signal input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew signal input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew signal input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew signal input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew signal input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew signal input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew signal input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew signal input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew signal input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew signal input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew signal input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew signal input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew signal input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew signal input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew signal input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew signal input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew signal input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew signal input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew signal input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew signal input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew signal input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew signal input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew signal input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew signal input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew signal input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew signal input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew signal input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew signal input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew signal input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew signal input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew signal input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew signal input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew signal input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew signal input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew signal input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew signal input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew signal input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew signal input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew signal input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew signal input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew signal input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew signal input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew signal input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew signal input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew signal input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew signal input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew signal input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew signal input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew signal input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew signal input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew signal input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew signal input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew signal input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew signal input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew signal input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew signal input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew signal input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew signal input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew signal input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew signal input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew signal input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew signal input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew signal input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew signal input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew signal input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew signal input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew signal input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew signal input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew signal input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew signal input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew signal input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew signal input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew signal input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew signal input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew signal input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew signal input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew signal input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew signal input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew signal input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew signal input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew signal input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew signal input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew signal input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew signal input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew signal input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew signal input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew signal input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew signal input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew signal input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew signal input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew signal input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew signal input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew signal input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew signal input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew signal input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew signal input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew signal input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew signal input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew signal input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew signal input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew signal input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew signal input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew signal input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew signal input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew signal input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew signal input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew signal input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew signal input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew signal input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew signal input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew signal input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew signal input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew signal input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew signal input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew signal input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew signal input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew signal input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew signal input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew signal input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew signal input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew signal input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew signal input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew signal input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew signal input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew signal input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew signal input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew signal input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew signal input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew signal input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew signal input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew signal input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew signal input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew signal input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew signal input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew signal input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew signal input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew signal input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew signal input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew signal input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew signal input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew signal input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew signal input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew signal input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew signal input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew signal input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew signal input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew signal input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew signal input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew signal input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew signal input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew signal input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew signal input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew signal input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew signal input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew signal tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew signal tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew signal tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew signal tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew signal tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew signal tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew signal tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew signal tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew signal tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew signal tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew signal tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew signal tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew signal tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew signal tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew signal tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew signal tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew signal tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew signal tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew signal tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew signal tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew signal tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew signal tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew signal tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew signal tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew signal tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew signal tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew signal tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew signal tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew signal tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew signal tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew signal tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew signal tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew signal input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew signal input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew signal input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew signal input
rlabel metal4 s 576804 -1864 577404 705800 6 vccd1
port 636 nsew power bidirectional
rlabel metal4 s 540804 -1864 541404 705800 6 vccd1.extra1
port 637 nsew power bidirectional
rlabel metal4 s 504804 -1864 505404 705800 6 vccd1.extra2
port 638 nsew power bidirectional
rlabel metal4 s 468804 -1864 469404 705800 6 vccd1.extra3
port 639 nsew power bidirectional
rlabel metal4 s 432804 -1864 433404 705800 6 vccd1.extra4
port 640 nsew power bidirectional
rlabel metal4 s 396804 -1864 397404 705800 6 vccd1.extra5
port 641 nsew power bidirectional
rlabel metal4 s 360804 -1864 361404 705800 6 vccd1.extra6
port 642 nsew power bidirectional
rlabel metal4 s 324804 -1864 325404 705800 6 vccd1.extra7
port 643 nsew power bidirectional
rlabel metal4 s 288804 -1864 289404 705800 6 vccd1.extra8
port 644 nsew power bidirectional
rlabel metal4 s 252804 267005 253404 705799 6 vccd1.extra9
port 645 nsew power bidirectional
rlabel metal4 s 216804 267005 217404 705799 6 vccd1.extra10
port 646 nsew power bidirectional
rlabel metal4 s 180804 267005 181404 705799 6 vccd1.extra11
port 647 nsew power bidirectional
rlabel metal4 s 144804 267005 145404 705799 6 vccd1.extra12
port 648 nsew power bidirectional
rlabel metal4 s 108804 267005 109404 705799 6 vccd1.extra13
port 649 nsew power bidirectional
rlabel metal4 s 72804 267005 73404 705799 6 vccd1.extra14
port 650 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 705800 6 vccd1.extra15
port 651 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 705800 6 vccd1.extra16
port 652 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1.extra17
port 653 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1.extra18
port 654 nsew power bidirectional
rlabel metal4 s 252804 -1864 253404 41200 6 vccd1.extra19
port 655 nsew power bidirectional
rlabel metal4 s 216804 -1864 217404 41200 6 vccd1.extra20
port 656 nsew power bidirectional
rlabel metal4 s 180804 -1864 181404 41200 6 vccd1.extra21
port 657 nsew power bidirectional
rlabel metal4 s 144804 -1864 145404 41200 6 vccd1.extra22
port 658 nsew power bidirectional
rlabel metal4 s 108804 -1864 109404 41200 6 vccd1.extra23
port 659 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 41200 6 vccd1.extra24
port 660 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1.extra25
port 661 nsew power bidirectional
rlabel metal5 s -2936 685876 586860 686476 6 vccd1.extra26
port 662 nsew power bidirectional
rlabel metal5 s -2936 649876 586860 650476 6 vccd1.extra27
port 663 nsew power bidirectional
rlabel metal5 s -2936 613876 586860 614476 6 vccd1.extra28
port 664 nsew power bidirectional
rlabel metal5 s -2936 577876 586860 578476 6 vccd1.extra29
port 665 nsew power bidirectional
rlabel metal5 s -2936 541876 586860 542476 6 vccd1.extra30
port 666 nsew power bidirectional
rlabel metal5 s -2936 505876 586860 506476 6 vccd1.extra31
port 667 nsew power bidirectional
rlabel metal5 s -2936 469876 586860 470476 6 vccd1.extra32
port 668 nsew power bidirectional
rlabel metal5 s -2936 433876 586860 434476 6 vccd1.extra33
port 669 nsew power bidirectional
rlabel metal5 s -2936 397876 586860 398476 6 vccd1.extra34
port 670 nsew power bidirectional
rlabel metal5 s -2936 361876 586860 362476 6 vccd1.extra35
port 671 nsew power bidirectional
rlabel metal5 s -2936 325876 586860 326476 6 vccd1.extra36
port 672 nsew power bidirectional
rlabel metal5 s -2936 289876 586860 290476 6 vccd1.extra37
port 673 nsew power bidirectional
rlabel metal5 s -2936 253876 586860 254476 6 vccd1.extra38
port 674 nsew power bidirectional
rlabel metal5 s -2936 217876 586860 218476 6 vccd1.extra39
port 675 nsew power bidirectional
rlabel metal5 s -2936 181876 586860 182476 6 vccd1.extra40
port 676 nsew power bidirectional
rlabel metal5 s -2936 145876 586860 146476 6 vccd1.extra41
port 677 nsew power bidirectional
rlabel metal5 s -2936 109876 586860 110476 6 vccd1.extra42
port 678 nsew power bidirectional
rlabel metal5 s -2936 73876 586860 74476 6 vccd1.extra43
port 679 nsew power bidirectional
rlabel metal5 s -2936 37876 586860 38476 6 vccd1.extra44
port 680 nsew power bidirectional
rlabel metal5 s -2936 1876 586860 2476 6 vccd1.extra45
port 681 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1.extra46
port 682 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 683 nsew ground bidirectional
rlabel metal4 s 558804 -1864 559404 705800 6 vssd1.extra1
port 684 nsew ground bidirectional
rlabel metal4 s 522804 -1864 523404 705800 6 vssd1.extra2
port 685 nsew ground bidirectional
rlabel metal4 s 486804 -1864 487404 705800 6 vssd1.extra3
port 686 nsew ground bidirectional
rlabel metal4 s 450804 -1864 451404 705800 6 vssd1.extra4
port 687 nsew ground bidirectional
rlabel metal4 s 414804 -1864 415404 705800 6 vssd1.extra5
port 688 nsew ground bidirectional
rlabel metal4 s 378804 -1864 379404 705800 6 vssd1.extra6
port 689 nsew ground bidirectional
rlabel metal4 s 342804 -1864 343404 705800 6 vssd1.extra7
port 690 nsew ground bidirectional
rlabel metal4 s 306804 -1864 307404 705800 6 vssd1.extra8
port 691 nsew ground bidirectional
rlabel metal4 s 270804 267005 271404 705799 6 vssd1.extra9
port 692 nsew ground bidirectional
rlabel metal4 s 234804 267005 235404 705799 6 vssd1.extra10
port 693 nsew ground bidirectional
rlabel metal4 s 198804 267005 199404 705799 6 vssd1.extra11
port 694 nsew ground bidirectional
rlabel metal4 s 162804 267005 163404 705799 6 vssd1.extra12
port 695 nsew ground bidirectional
rlabel metal4 s 126804 267005 127404 705799 6 vssd1.extra13
port 696 nsew ground bidirectional
rlabel metal4 s 90804 267005 91404 705799 6 vssd1.extra14
port 697 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 705800 6 vssd1.extra15
port 698 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 705800 6 vssd1.extra16
port 699 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1.extra17
port 700 nsew ground bidirectional
rlabel metal4 s 270804 -1864 271404 41200 6 vssd1.extra18
port 701 nsew ground bidirectional
rlabel metal4 s 234804 -1864 235404 41200 6 vssd1.extra19
port 702 nsew ground bidirectional
rlabel metal4 s 198804 -1864 199404 41200 6 vssd1.extra20
port 703 nsew ground bidirectional
rlabel metal4 s 162804 -1864 163404 41200 6 vssd1.extra21
port 704 nsew ground bidirectional
rlabel metal4 s 126804 -1864 127404 41200 6 vssd1.extra22
port 705 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 41200 6 vssd1.extra23
port 706 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1.extra24
port 707 nsew ground bidirectional
rlabel metal5 s -2936 667876 586860 668476 6 vssd1.extra25
port 708 nsew ground bidirectional
rlabel metal5 s -2936 631876 586860 632476 6 vssd1.extra26
port 709 nsew ground bidirectional
rlabel metal5 s -2936 595876 586860 596476 6 vssd1.extra27
port 710 nsew ground bidirectional
rlabel metal5 s -2936 559876 586860 560476 6 vssd1.extra28
port 711 nsew ground bidirectional
rlabel metal5 s -2936 523876 586860 524476 6 vssd1.extra29
port 712 nsew ground bidirectional
rlabel metal5 s -2936 487876 586860 488476 6 vssd1.extra30
port 713 nsew ground bidirectional
rlabel metal5 s -2936 451876 586860 452476 6 vssd1.extra31
port 714 nsew ground bidirectional
rlabel metal5 s -2936 415876 586860 416476 6 vssd1.extra32
port 715 nsew ground bidirectional
rlabel metal5 s -2936 379876 586860 380476 6 vssd1.extra33
port 716 nsew ground bidirectional
rlabel metal5 s -2936 343876 586860 344476 6 vssd1.extra34
port 717 nsew ground bidirectional
rlabel metal5 s -2936 307876 586860 308476 6 vssd1.extra35
port 718 nsew ground bidirectional
rlabel metal5 s -2936 271876 586860 272476 6 vssd1.extra36
port 719 nsew ground bidirectional
rlabel metal5 s -2936 235876 586860 236476 6 vssd1.extra37
port 720 nsew ground bidirectional
rlabel metal5 s -2936 199876 586860 200476 6 vssd1.extra38
port 721 nsew ground bidirectional
rlabel metal5 s -2936 163876 586860 164476 6 vssd1.extra39
port 722 nsew ground bidirectional
rlabel metal5 s -2936 127876 586860 128476 6 vssd1.extra40
port 723 nsew ground bidirectional
rlabel metal5 s -2936 91876 586860 92476 6 vssd1.extra41
port 724 nsew ground bidirectional
rlabel metal5 s -2936 55876 586860 56476 6 vssd1.extra42
port 725 nsew ground bidirectional
rlabel metal5 s -2936 19876 586860 20476 6 vssd1.extra43
port 726 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1.extra44
port 727 nsew ground bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 728 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2.extra1
port 729 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2.extra2
port 730 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2.extra3
port 731 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 732 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2.extra1
port 733 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2.extra2
port 734 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2.extra3
port 735 nsew ground bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 736 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1.extra1
port 737 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1.extra2
port 738 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1.extra3
port 739 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 740 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1.extra1
port 741 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1.extra2
port 742 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1.extra3
port 743 nsew ground bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 744 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2.extra1
port 745 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2.extra2
port 746 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2.extra3
port 747 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 748 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2.extra1
port 749 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2.extra2
port 750 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2.extra3
port 751 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
