VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 279.750 503.780 280.070 503.840 ;
        RECT 296.770 503.780 297.090 503.840 ;
        RECT 279.750 503.640 297.090 503.780 ;
        RECT 279.750 503.580 280.070 503.640 ;
        RECT 296.770 503.580 297.090 503.640 ;
        RECT 279.750 89.660 280.070 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 279.750 89.520 2899.310 89.660 ;
        RECT 279.750 89.460 280.070 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 279.780 503.580 280.040 503.840 ;
        RECT 296.800 503.580 297.060 503.840 ;
        RECT 279.780 89.460 280.040 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 296.790 504.715 297.070 505.085 ;
        RECT 296.860 503.870 297.000 504.715 ;
        RECT 279.780 503.550 280.040 503.870 ;
        RECT 296.800 503.550 297.060 503.870 ;
        RECT 279.840 89.750 279.980 503.550 ;
        RECT 279.780 89.430 280.040 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 296.790 504.760 297.070 505.040 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 296.765 505.050 297.095 505.065 ;
        RECT 296.765 504.960 310.500 505.050 ;
        RECT 296.765 504.750 314.000 504.960 ;
        RECT 296.765 504.735 297.095 504.750 ;
        RECT 310.000 504.360 314.000 504.750 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1459.190 2429.200 1459.510 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 1459.190 2429.060 2901.150 2429.200 ;
        RECT 1459.190 2429.000 1459.510 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 1098.550 198.460 1098.870 198.520 ;
        RECT 1459.190 198.460 1459.510 198.520 ;
        RECT 1098.550 198.320 1459.510 198.460 ;
        RECT 1098.550 198.260 1098.870 198.320 ;
        RECT 1459.190 198.260 1459.510 198.320 ;
      LAYER via ;
        RECT 1459.220 2429.000 1459.480 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 1098.580 198.260 1098.840 198.520 ;
        RECT 1459.220 198.260 1459.480 198.520 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 1459.220 2428.970 1459.480 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 1098.530 216.000 1098.810 220.000 ;
        RECT 1098.640 198.550 1098.780 216.000 ;
        RECT 1459.280 198.550 1459.420 2428.970 ;
        RECT 1098.580 198.230 1098.840 198.550 ;
        RECT 1459.220 198.230 1459.480 198.550 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1248.510 2663.800 1248.830 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 1248.510 2663.660 2901.150 2663.800 ;
        RECT 1248.510 2663.600 1248.830 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
        RECT 1244.830 1338.480 1245.150 1338.540 ;
        RECT 1248.510 1338.480 1248.830 1338.540 ;
        RECT 1244.830 1338.340 1248.830 1338.480 ;
        RECT 1244.830 1338.280 1245.150 1338.340 ;
        RECT 1248.510 1338.280 1248.830 1338.340 ;
      LAYER via ;
        RECT 1248.540 2663.600 1248.800 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
        RECT 1244.860 1338.280 1245.120 1338.540 ;
        RECT 1248.540 1338.280 1248.800 1338.540 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 1248.540 2663.570 1248.800 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 1248.600 1338.570 1248.740 2663.570 ;
        RECT 1244.860 1338.250 1245.120 1338.570 ;
        RECT 1248.540 1338.250 1248.800 1338.570 ;
        RECT 1244.920 1325.025 1245.060 1338.250 ;
        RECT 1244.810 1321.025 1245.090 1325.025 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1645.490 2898.400 1645.810 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 1645.490 2898.260 2901.150 2898.400 ;
        RECT 1645.490 2898.200 1645.810 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 1325.790 199.820 1326.110 199.880 ;
        RECT 1645.490 199.820 1645.810 199.880 ;
        RECT 1325.790 199.680 1645.810 199.820 ;
        RECT 1325.790 199.620 1326.110 199.680 ;
        RECT 1645.490 199.620 1645.810 199.680 ;
      LAYER via ;
        RECT 1645.520 2898.200 1645.780 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 1325.820 199.620 1326.080 199.880 ;
        RECT 1645.520 199.620 1645.780 199.880 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 1645.520 2898.170 1645.780 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 1325.770 216.000 1326.050 220.000 ;
        RECT 1325.880 199.910 1326.020 216.000 ;
        RECT 1645.580 199.910 1645.720 2898.170 ;
        RECT 1325.820 199.590 1326.080 199.910 ;
        RECT 1645.520 199.590 1645.780 199.910 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1424.690 3133.000 1425.010 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 1424.690 3132.860 2901.150 3133.000 ;
        RECT 1424.690 3132.800 1425.010 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
        RECT 371.750 198.800 372.070 198.860 ;
        RECT 1424.690 198.800 1425.010 198.860 ;
        RECT 371.750 198.660 1425.010 198.800 ;
        RECT 371.750 198.600 372.070 198.660 ;
        RECT 1424.690 198.600 1425.010 198.660 ;
      LAYER via ;
        RECT 1424.720 3132.800 1424.980 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
        RECT 371.780 198.600 372.040 198.860 ;
        RECT 1424.720 198.600 1424.980 198.860 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 1424.720 3132.770 1424.980 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 371.730 216.000 372.010 220.000 ;
        RECT 371.840 198.890 371.980 216.000 ;
        RECT 1424.780 198.890 1424.920 3132.770 ;
        RECT 371.780 198.570 372.040 198.890 ;
        RECT 1424.720 198.570 1424.980 198.890 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 303.210 3367.600 303.530 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 303.210 3367.460 2901.150 3367.600 ;
        RECT 303.210 3367.400 303.530 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 303.240 3367.400 303.500 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 303.240 3367.370 303.500 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 303.300 864.125 303.440 3367.370 ;
        RECT 303.230 863.755 303.510 864.125 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 303.230 863.800 303.510 864.080 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 303.205 864.090 303.535 864.105 ;
        RECT 303.205 864.000 310.500 864.090 ;
        RECT 303.205 863.790 314.000 864.000 ;
        RECT 303.205 863.775 303.535 863.790 ;
        RECT 310.000 863.400 314.000 863.790 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2666.690 3501.560 2667.010 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 2666.690 3501.420 2798.570 3501.560 ;
        RECT 2666.690 3501.360 2667.010 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
        RECT 475.710 200.160 476.030 200.220 ;
        RECT 2666.690 200.160 2667.010 200.220 ;
        RECT 475.710 200.020 2667.010 200.160 ;
        RECT 475.710 199.960 476.030 200.020 ;
        RECT 2666.690 199.960 2667.010 200.020 ;
      LAYER via ;
        RECT 2666.720 3501.360 2666.980 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
        RECT 475.740 199.960 476.000 200.220 ;
        RECT 2666.720 199.960 2666.980 200.220 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 2666.720 3501.330 2666.980 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 475.690 216.000 475.970 220.000 ;
        RECT 475.800 200.250 475.940 216.000 ;
        RECT 2666.780 200.250 2666.920 3501.330 ;
        RECT 475.740 199.930 476.000 200.250 ;
        RECT 2666.720 199.930 2666.980 200.250 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
        RECT 2471.265 2753.065 2471.435 2767.175 ;
        RECT 2471.265 1787.465 2471.435 1801.235 ;
        RECT 2470.345 1690.565 2470.515 1738.675 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
        RECT 2471.265 2767.005 2471.435 2767.175 ;
        RECT 2471.265 1801.065 2471.435 1801.235 ;
        RECT 2470.345 1738.505 2470.515 1738.675 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 3077.580 2470.590 3077.640 ;
        RECT 2471.190 3077.580 2471.510 3077.640 ;
        RECT 2470.270 3077.440 2471.510 3077.580 ;
        RECT 2470.270 3077.380 2470.590 3077.440 ;
        RECT 2471.190 3077.380 2471.510 3077.440 ;
        RECT 2470.270 2981.020 2470.590 2981.080 ;
        RECT 2471.190 2981.020 2471.510 2981.080 ;
        RECT 2470.270 2980.880 2471.510 2981.020 ;
        RECT 2470.270 2980.820 2470.590 2980.880 ;
        RECT 2471.190 2980.820 2471.510 2980.880 ;
        RECT 2469.350 2946.340 2469.670 2946.400 ;
        RECT 2470.730 2946.340 2471.050 2946.400 ;
        RECT 2469.350 2946.200 2471.050 2946.340 ;
        RECT 2469.350 2946.140 2469.670 2946.200 ;
        RECT 2470.730 2946.140 2471.050 2946.200 ;
        RECT 2471.190 2767.160 2471.510 2767.220 ;
        RECT 2470.995 2767.020 2471.510 2767.160 ;
        RECT 2471.190 2766.960 2471.510 2767.020 ;
        RECT 2471.190 2753.220 2471.510 2753.280 ;
        RECT 2470.995 2753.080 2471.510 2753.220 ;
        RECT 2471.190 2753.020 2471.510 2753.080 ;
        RECT 2471.190 2719.020 2471.510 2719.280 ;
        RECT 2471.280 2718.880 2471.420 2719.020 ;
        RECT 2471.650 2718.880 2471.970 2718.940 ;
        RECT 2471.280 2718.740 2471.970 2718.880 ;
        RECT 2471.650 2718.680 2471.970 2718.740 ;
        RECT 2470.730 2656.660 2471.050 2656.720 ;
        RECT 2472.110 2656.660 2472.430 2656.720 ;
        RECT 2470.730 2656.520 2472.430 2656.660 ;
        RECT 2470.730 2656.460 2471.050 2656.520 ;
        RECT 2472.110 2656.460 2472.430 2656.520 ;
        RECT 2472.110 2622.660 2472.430 2622.720 ;
        RECT 2471.740 2622.520 2472.430 2622.660 ;
        RECT 2471.740 2622.040 2471.880 2622.520 ;
        RECT 2472.110 2622.460 2472.430 2622.520 ;
        RECT 2471.650 2621.780 2471.970 2622.040 ;
        RECT 2470.730 2560.100 2471.050 2560.160 ;
        RECT 2472.110 2560.100 2472.430 2560.160 ;
        RECT 2470.730 2559.960 2472.430 2560.100 ;
        RECT 2470.730 2559.900 2471.050 2559.960 ;
        RECT 2472.110 2559.900 2472.430 2559.960 ;
        RECT 2471.190 2511.820 2471.510 2511.880 ;
        RECT 2472.110 2511.820 2472.430 2511.880 ;
        RECT 2471.190 2511.680 2472.430 2511.820 ;
        RECT 2471.190 2511.620 2471.510 2511.680 ;
        RECT 2472.110 2511.620 2472.430 2511.680 ;
        RECT 2470.270 2401.320 2470.590 2401.380 ;
        RECT 2471.190 2401.320 2471.510 2401.380 ;
        RECT 2470.270 2401.180 2471.510 2401.320 ;
        RECT 2470.270 2401.120 2470.590 2401.180 ;
        RECT 2471.190 2401.120 2471.510 2401.180 ;
        RECT 2470.270 2304.760 2470.590 2304.820 ;
        RECT 2471.190 2304.760 2471.510 2304.820 ;
        RECT 2470.270 2304.620 2471.510 2304.760 ;
        RECT 2470.270 2304.560 2470.590 2304.620 ;
        RECT 2471.190 2304.560 2471.510 2304.620 ;
        RECT 2470.270 2208.200 2470.590 2208.260 ;
        RECT 2471.190 2208.200 2471.510 2208.260 ;
        RECT 2470.270 2208.060 2471.510 2208.200 ;
        RECT 2470.270 2208.000 2470.590 2208.060 ;
        RECT 2471.190 2208.000 2471.510 2208.060 ;
        RECT 2470.270 2111.640 2470.590 2111.700 ;
        RECT 2471.190 2111.640 2471.510 2111.700 ;
        RECT 2470.270 2111.500 2471.510 2111.640 ;
        RECT 2470.270 2111.440 2470.590 2111.500 ;
        RECT 2471.190 2111.440 2471.510 2111.500 ;
        RECT 2470.270 2015.080 2470.590 2015.140 ;
        RECT 2471.190 2015.080 2471.510 2015.140 ;
        RECT 2470.270 2014.940 2471.510 2015.080 ;
        RECT 2470.270 2014.880 2470.590 2014.940 ;
        RECT 2471.190 2014.880 2471.510 2014.940 ;
        RECT 2470.270 1918.520 2470.590 1918.580 ;
        RECT 2471.190 1918.520 2471.510 1918.580 ;
        RECT 2470.270 1918.380 2471.510 1918.520 ;
        RECT 2470.270 1918.320 2470.590 1918.380 ;
        RECT 2471.190 1918.320 2471.510 1918.380 ;
        RECT 2471.190 1801.220 2471.510 1801.280 ;
        RECT 2470.995 1801.080 2471.510 1801.220 ;
        RECT 2471.190 1801.020 2471.510 1801.080 ;
        RECT 2471.190 1787.620 2471.510 1787.680 ;
        RECT 2470.995 1787.480 2471.510 1787.620 ;
        RECT 2471.190 1787.420 2471.510 1787.480 ;
        RECT 2470.270 1738.660 2470.590 1738.720 ;
        RECT 2470.075 1738.520 2470.590 1738.660 ;
        RECT 2470.270 1738.460 2470.590 1738.520 ;
        RECT 2470.285 1690.720 2470.575 1690.765 ;
        RECT 2470.730 1690.720 2471.050 1690.780 ;
        RECT 2470.285 1690.580 2471.050 1690.720 ;
        RECT 2470.285 1690.535 2470.575 1690.580 ;
        RECT 2470.730 1690.520 2471.050 1690.580 ;
        RECT 2470.270 1628.500 2470.590 1628.560 ;
        RECT 2471.190 1628.500 2471.510 1628.560 ;
        RECT 2470.270 1628.360 2471.510 1628.500 ;
        RECT 2470.270 1628.300 2470.590 1628.360 ;
        RECT 2471.190 1628.300 2471.510 1628.360 ;
        RECT 2470.270 1531.940 2470.590 1532.000 ;
        RECT 2471.190 1531.940 2471.510 1532.000 ;
        RECT 2470.270 1531.800 2471.510 1531.940 ;
        RECT 2470.270 1531.740 2470.590 1531.800 ;
        RECT 2471.190 1531.740 2471.510 1531.800 ;
        RECT 2470.270 1435.380 2470.590 1435.440 ;
        RECT 2471.190 1435.380 2471.510 1435.440 ;
        RECT 2470.270 1435.240 2471.510 1435.380 ;
        RECT 2470.270 1435.180 2470.590 1435.240 ;
        RECT 2471.190 1435.180 2471.510 1435.240 ;
        RECT 1432.510 1410.900 1432.830 1410.960 ;
        RECT 2470.270 1410.900 2470.590 1410.960 ;
        RECT 1432.510 1410.760 2470.590 1410.900 ;
        RECT 1432.510 1410.700 1432.830 1410.760 ;
        RECT 2470.270 1410.700 2470.590 1410.760 ;
        RECT 1420.550 1142.980 1420.870 1143.040 ;
        RECT 1432.510 1142.980 1432.830 1143.040 ;
        RECT 1420.550 1142.840 1432.830 1142.980 ;
        RECT 1420.550 1142.780 1420.870 1142.840 ;
        RECT 1432.510 1142.780 1432.830 1142.840 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 3077.380 2470.560 3077.640 ;
        RECT 2471.220 3077.380 2471.480 3077.640 ;
        RECT 2470.300 2980.820 2470.560 2981.080 ;
        RECT 2471.220 2980.820 2471.480 2981.080 ;
        RECT 2469.380 2946.140 2469.640 2946.400 ;
        RECT 2470.760 2946.140 2471.020 2946.400 ;
        RECT 2471.220 2766.960 2471.480 2767.220 ;
        RECT 2471.220 2753.020 2471.480 2753.280 ;
        RECT 2471.220 2719.020 2471.480 2719.280 ;
        RECT 2471.680 2718.680 2471.940 2718.940 ;
        RECT 2470.760 2656.460 2471.020 2656.720 ;
        RECT 2472.140 2656.460 2472.400 2656.720 ;
        RECT 2472.140 2622.460 2472.400 2622.720 ;
        RECT 2471.680 2621.780 2471.940 2622.040 ;
        RECT 2470.760 2559.900 2471.020 2560.160 ;
        RECT 2472.140 2559.900 2472.400 2560.160 ;
        RECT 2471.220 2511.620 2471.480 2511.880 ;
        RECT 2472.140 2511.620 2472.400 2511.880 ;
        RECT 2470.300 2401.120 2470.560 2401.380 ;
        RECT 2471.220 2401.120 2471.480 2401.380 ;
        RECT 2470.300 2304.560 2470.560 2304.820 ;
        RECT 2471.220 2304.560 2471.480 2304.820 ;
        RECT 2470.300 2208.000 2470.560 2208.260 ;
        RECT 2471.220 2208.000 2471.480 2208.260 ;
        RECT 2470.300 2111.440 2470.560 2111.700 ;
        RECT 2471.220 2111.440 2471.480 2111.700 ;
        RECT 2470.300 2014.880 2470.560 2015.140 ;
        RECT 2471.220 2014.880 2471.480 2015.140 ;
        RECT 2470.300 1918.320 2470.560 1918.580 ;
        RECT 2471.220 1918.320 2471.480 1918.580 ;
        RECT 2471.220 1801.020 2471.480 1801.280 ;
        RECT 2471.220 1787.420 2471.480 1787.680 ;
        RECT 2470.300 1738.460 2470.560 1738.720 ;
        RECT 2470.760 1690.520 2471.020 1690.780 ;
        RECT 2470.300 1628.300 2470.560 1628.560 ;
        RECT 2471.220 1628.300 2471.480 1628.560 ;
        RECT 2470.300 1531.740 2470.560 1532.000 ;
        RECT 2471.220 1531.740 2471.480 1532.000 ;
        RECT 2470.300 1435.180 2470.560 1435.440 ;
        RECT 2471.220 1435.180 2471.480 1435.440 ;
        RECT 1432.540 1410.700 1432.800 1410.960 ;
        RECT 2470.300 1410.700 2470.560 1410.960 ;
        RECT 1420.580 1142.780 1420.840 1143.040 ;
        RECT 1432.540 1142.780 1432.800 1143.040 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3430.445 2474.640 3517.230 ;
        RECT 2474.430 3430.075 2474.710 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3298.410 2470.960 3332.690 ;
        RECT 2470.820 3298.270 2471.420 3298.410 ;
        RECT 2471.280 3270.790 2471.420 3298.270 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3222.250 2470.500 3270.470 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 3077.670 2471.420 3125.550 ;
        RECT 2470.300 3077.350 2470.560 3077.670 ;
        RECT 2471.220 3077.350 2471.480 3077.670 ;
        RECT 2470.360 3029.130 2470.500 3077.350 ;
        RECT 2470.360 3028.990 2471.420 3029.130 ;
        RECT 2471.280 2981.110 2471.420 3028.990 ;
        RECT 2470.300 2980.850 2470.560 2981.110 ;
        RECT 2470.300 2980.790 2470.960 2980.850 ;
        RECT 2471.220 2980.790 2471.480 2981.110 ;
        RECT 2470.360 2980.710 2470.960 2980.790 ;
        RECT 2470.820 2980.170 2470.960 2980.710 ;
        RECT 2470.820 2980.030 2471.420 2980.170 ;
        RECT 2471.280 2959.770 2471.420 2980.030 ;
        RECT 2470.820 2959.630 2471.420 2959.770 ;
        RECT 2470.820 2946.430 2470.960 2959.630 ;
        RECT 2469.380 2946.110 2469.640 2946.430 ;
        RECT 2470.760 2946.110 2471.020 2946.430 ;
        RECT 2469.440 2898.685 2469.580 2946.110 ;
        RECT 2469.370 2898.315 2469.650 2898.685 ;
        RECT 2470.290 2898.315 2470.570 2898.685 ;
        RECT 2470.360 2863.210 2470.500 2898.315 ;
        RECT 2470.360 2863.070 2470.960 2863.210 ;
        RECT 2470.820 2815.610 2470.960 2863.070 ;
        RECT 2470.820 2815.470 2471.420 2815.610 ;
        RECT 2471.280 2767.250 2471.420 2815.470 ;
        RECT 2471.220 2766.930 2471.480 2767.250 ;
        RECT 2471.220 2752.990 2471.480 2753.310 ;
        RECT 2471.280 2719.310 2471.420 2752.990 ;
        RECT 2471.220 2718.990 2471.480 2719.310 ;
        RECT 2471.680 2718.650 2471.940 2718.970 ;
        RECT 2471.740 2704.885 2471.880 2718.650 ;
        RECT 2470.750 2704.515 2471.030 2704.885 ;
        RECT 2471.670 2704.515 2471.950 2704.885 ;
        RECT 2470.820 2656.750 2470.960 2704.515 ;
        RECT 2470.760 2656.430 2471.020 2656.750 ;
        RECT 2472.140 2656.430 2472.400 2656.750 ;
        RECT 2472.200 2622.750 2472.340 2656.430 ;
        RECT 2472.140 2622.430 2472.400 2622.750 ;
        RECT 2471.680 2621.750 2471.940 2622.070 ;
        RECT 2471.740 2608.325 2471.880 2621.750 ;
        RECT 2470.750 2607.955 2471.030 2608.325 ;
        RECT 2471.670 2607.955 2471.950 2608.325 ;
        RECT 2470.820 2560.190 2470.960 2607.955 ;
        RECT 2470.760 2559.870 2471.020 2560.190 ;
        RECT 2472.140 2559.870 2472.400 2560.190 ;
        RECT 2472.200 2511.910 2472.340 2559.870 ;
        RECT 2471.220 2511.765 2471.480 2511.910 ;
        RECT 2469.830 2511.395 2470.110 2511.765 ;
        RECT 2471.210 2511.395 2471.490 2511.765 ;
        RECT 2472.140 2511.590 2472.400 2511.910 ;
        RECT 2469.900 2463.485 2470.040 2511.395 ;
        RECT 2469.830 2463.115 2470.110 2463.485 ;
        RECT 2470.750 2463.115 2471.030 2463.485 ;
        RECT 2470.820 2449.770 2470.960 2463.115 ;
        RECT 2470.820 2449.630 2471.420 2449.770 ;
        RECT 2471.280 2401.410 2471.420 2449.630 ;
        RECT 2470.300 2401.090 2470.560 2401.410 ;
        RECT 2471.220 2401.090 2471.480 2401.410 ;
        RECT 2470.360 2400.810 2470.500 2401.090 ;
        RECT 2470.360 2400.670 2470.960 2400.810 ;
        RECT 2470.820 2353.210 2470.960 2400.670 ;
        RECT 2470.820 2353.070 2471.420 2353.210 ;
        RECT 2471.280 2304.850 2471.420 2353.070 ;
        RECT 2470.300 2304.530 2470.560 2304.850 ;
        RECT 2471.220 2304.530 2471.480 2304.850 ;
        RECT 2470.360 2304.250 2470.500 2304.530 ;
        RECT 2470.360 2304.110 2470.960 2304.250 ;
        RECT 2470.820 2256.650 2470.960 2304.110 ;
        RECT 2470.820 2256.510 2471.420 2256.650 ;
        RECT 2471.280 2208.290 2471.420 2256.510 ;
        RECT 2470.300 2207.970 2470.560 2208.290 ;
        RECT 2471.220 2207.970 2471.480 2208.290 ;
        RECT 2470.360 2207.690 2470.500 2207.970 ;
        RECT 2470.360 2207.550 2470.960 2207.690 ;
        RECT 2470.820 2160.090 2470.960 2207.550 ;
        RECT 2470.820 2159.950 2471.420 2160.090 ;
        RECT 2471.280 2111.730 2471.420 2159.950 ;
        RECT 2470.300 2111.410 2470.560 2111.730 ;
        RECT 2471.220 2111.410 2471.480 2111.730 ;
        RECT 2470.360 2111.130 2470.500 2111.410 ;
        RECT 2470.360 2110.990 2470.960 2111.130 ;
        RECT 2470.820 2063.530 2470.960 2110.990 ;
        RECT 2470.820 2063.390 2471.420 2063.530 ;
        RECT 2471.280 2015.170 2471.420 2063.390 ;
        RECT 2470.300 2014.850 2470.560 2015.170 ;
        RECT 2471.220 2014.850 2471.480 2015.170 ;
        RECT 2470.360 2014.570 2470.500 2014.850 ;
        RECT 2470.360 2014.430 2470.960 2014.570 ;
        RECT 2470.820 1966.970 2470.960 2014.430 ;
        RECT 2470.820 1966.830 2471.420 1966.970 ;
        RECT 2471.280 1918.610 2471.420 1966.830 ;
        RECT 2470.300 1918.290 2470.560 1918.610 ;
        RECT 2471.220 1918.290 2471.480 1918.610 ;
        RECT 2470.360 1918.010 2470.500 1918.290 ;
        RECT 2470.360 1917.870 2470.960 1918.010 ;
        RECT 2470.820 1870.410 2470.960 1917.870 ;
        RECT 2470.820 1870.270 2471.420 1870.410 ;
        RECT 2471.280 1801.310 2471.420 1870.270 ;
        RECT 2471.220 1800.990 2471.480 1801.310 ;
        RECT 2471.220 1787.390 2471.480 1787.710 ;
        RECT 2471.280 1752.770 2471.420 1787.390 ;
        RECT 2470.360 1752.630 2471.420 1752.770 ;
        RECT 2470.360 1738.750 2470.500 1752.630 ;
        RECT 2470.300 1738.430 2470.560 1738.750 ;
        RECT 2470.760 1690.490 2471.020 1690.810 ;
        RECT 2470.820 1656.210 2470.960 1690.490 ;
        RECT 2470.820 1656.070 2471.420 1656.210 ;
        RECT 2471.280 1628.590 2471.420 1656.070 ;
        RECT 2470.300 1628.270 2470.560 1628.590 ;
        RECT 2471.220 1628.270 2471.480 1628.590 ;
        RECT 2470.360 1580.050 2470.500 1628.270 ;
        RECT 2470.360 1579.910 2471.420 1580.050 ;
        RECT 2471.280 1532.030 2471.420 1579.910 ;
        RECT 2470.300 1531.710 2470.560 1532.030 ;
        RECT 2471.220 1531.710 2471.480 1532.030 ;
        RECT 2470.360 1483.490 2470.500 1531.710 ;
        RECT 2470.360 1483.350 2471.420 1483.490 ;
        RECT 2471.280 1435.470 2471.420 1483.350 ;
        RECT 2470.300 1435.150 2470.560 1435.470 ;
        RECT 2471.220 1435.150 2471.480 1435.470 ;
        RECT 2470.360 1410.990 2470.500 1435.150 ;
        RECT 1432.540 1410.670 1432.800 1410.990 ;
        RECT 2470.300 1410.670 2470.560 1410.990 ;
        RECT 1432.600 1143.070 1432.740 1410.670 ;
        RECT 1420.580 1142.750 1420.840 1143.070 ;
        RECT 1432.540 1142.750 1432.800 1143.070 ;
        RECT 1420.640 1141.565 1420.780 1142.750 ;
        RECT 1420.570 1141.195 1420.850 1141.565 ;
      LAYER via2 ;
        RECT 2474.430 3430.120 2474.710 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
        RECT 2469.370 2898.360 2469.650 2898.640 ;
        RECT 2470.290 2898.360 2470.570 2898.640 ;
        RECT 2470.750 2704.560 2471.030 2704.840 ;
        RECT 2471.670 2704.560 2471.950 2704.840 ;
        RECT 2470.750 2608.000 2471.030 2608.280 ;
        RECT 2471.670 2608.000 2471.950 2608.280 ;
        RECT 2469.830 2511.440 2470.110 2511.720 ;
        RECT 2471.210 2511.440 2471.490 2511.720 ;
        RECT 2469.830 2463.160 2470.110 2463.440 ;
        RECT 2470.750 2463.160 2471.030 2463.440 ;
        RECT 1420.570 1141.240 1420.850 1141.520 ;
      LAYER met3 ;
        RECT 2474.405 3430.410 2474.735 3430.425 ;
        RECT 2470.510 3430.110 2474.735 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.405 3430.095 2474.735 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
        RECT 2469.345 2898.650 2469.675 2898.665 ;
        RECT 2470.265 2898.650 2470.595 2898.665 ;
        RECT 2469.345 2898.350 2470.595 2898.650 ;
        RECT 2469.345 2898.335 2469.675 2898.350 ;
        RECT 2470.265 2898.335 2470.595 2898.350 ;
        RECT 2470.725 2704.850 2471.055 2704.865 ;
        RECT 2471.645 2704.850 2471.975 2704.865 ;
        RECT 2470.725 2704.550 2471.975 2704.850 ;
        RECT 2470.725 2704.535 2471.055 2704.550 ;
        RECT 2471.645 2704.535 2471.975 2704.550 ;
        RECT 2470.725 2608.290 2471.055 2608.305 ;
        RECT 2471.645 2608.290 2471.975 2608.305 ;
        RECT 2470.725 2607.990 2471.975 2608.290 ;
        RECT 2470.725 2607.975 2471.055 2607.990 ;
        RECT 2471.645 2607.975 2471.975 2607.990 ;
        RECT 2469.805 2511.730 2470.135 2511.745 ;
        RECT 2471.185 2511.730 2471.515 2511.745 ;
        RECT 2469.805 2511.430 2471.515 2511.730 ;
        RECT 2469.805 2511.415 2470.135 2511.430 ;
        RECT 2471.185 2511.415 2471.515 2511.430 ;
        RECT 2469.805 2463.450 2470.135 2463.465 ;
        RECT 2470.725 2463.450 2471.055 2463.465 ;
        RECT 2469.805 2463.150 2471.055 2463.450 ;
        RECT 2469.805 2463.135 2470.135 2463.150 ;
        RECT 2470.725 2463.135 2471.055 2463.150 ;
        RECT 1420.545 1141.530 1420.875 1141.545 ;
        RECT 1408.060 1141.440 1420.875 1141.530 ;
        RECT 1404.305 1141.230 1420.875 1141.440 ;
        RECT 1404.305 1140.840 1408.305 1141.230 ;
        RECT 1420.545 1141.215 1420.875 1141.230 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3422.355 ;
        RECT 2146.965 3008.405 2147.135 3042.915 ;
        RECT 2147.885 2946.525 2148.055 2994.635 ;
        RECT 2146.505 2753.065 2146.675 2801.175 ;
        RECT 2146.965 2428.705 2147.135 2463.215 ;
        RECT 2146.965 2331.805 2147.135 2366.655 ;
        RECT 2146.505 1993.845 2146.675 2028.355 ;
        RECT 2147.885 1766.725 2148.055 1787.635 ;
        RECT 2148.345 1703.825 2148.515 1766.215 ;
        RECT 2147.425 1400.885 2147.595 1448.995 ;
        RECT 2146.965 1317.585 2147.135 1352.435 ;
        RECT 2147.885 1269.645 2148.055 1304.155 ;
        RECT 2146.505 1110.865 2146.675 1158.975 ;
        RECT 2147.425 966.365 2147.595 1014.135 ;
        RECT 2147.425 869.805 2147.595 917.575 ;
        RECT 2146.965 786.505 2147.135 821.015 ;
        RECT 2146.965 689.605 2147.135 724.455 ;
        RECT 2146.505 579.785 2146.675 627.895 ;
      LAYER mcon ;
        RECT 2147.885 3422.185 2148.055 3422.355 ;
        RECT 2146.965 3042.745 2147.135 3042.915 ;
        RECT 2147.885 2994.465 2148.055 2994.635 ;
        RECT 2146.505 2801.005 2146.675 2801.175 ;
        RECT 2146.965 2463.045 2147.135 2463.215 ;
        RECT 2146.965 2366.485 2147.135 2366.655 ;
        RECT 2146.505 2028.185 2146.675 2028.355 ;
        RECT 2147.885 1787.465 2148.055 1787.635 ;
        RECT 2148.345 1766.045 2148.515 1766.215 ;
        RECT 2147.425 1448.825 2147.595 1448.995 ;
        RECT 2146.965 1352.265 2147.135 1352.435 ;
        RECT 2147.885 1303.985 2148.055 1304.155 ;
        RECT 2146.505 1158.805 2146.675 1158.975 ;
        RECT 2147.425 1013.965 2147.595 1014.135 ;
        RECT 2147.425 917.405 2147.595 917.575 ;
        RECT 2146.965 820.845 2147.135 821.015 ;
        RECT 2146.965 724.285 2147.135 724.455 ;
        RECT 2146.505 627.725 2146.675 627.895 ;
      LAYER met1 ;
        RECT 2146.890 3443.080 2147.210 3443.140 ;
        RECT 2149.190 3443.080 2149.510 3443.140 ;
        RECT 2146.890 3442.940 2149.510 3443.080 ;
        RECT 2146.890 3442.880 2147.210 3442.940 ;
        RECT 2149.190 3442.880 2149.510 3442.940 ;
        RECT 2146.430 3422.340 2146.750 3422.400 ;
        RECT 2147.825 3422.340 2148.115 3422.385 ;
        RECT 2146.430 3422.200 2148.115 3422.340 ;
        RECT 2146.430 3422.140 2146.750 3422.200 ;
        RECT 2147.825 3422.155 2148.115 3422.200 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2146.430 3056.840 2146.750 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2146.430 3056.700 2147.670 3056.840 ;
        RECT 2146.430 3056.640 2146.750 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 2146.890 3042.900 2147.210 3042.960 ;
        RECT 2146.695 3042.760 2147.210 3042.900 ;
        RECT 2146.890 3042.700 2147.210 3042.760 ;
        RECT 2146.905 3008.560 2147.195 3008.605 ;
        RECT 2147.810 3008.560 2148.130 3008.620 ;
        RECT 2146.905 3008.420 2148.130 3008.560 ;
        RECT 2146.905 3008.375 2147.195 3008.420 ;
        RECT 2147.810 3008.360 2148.130 3008.420 ;
        RECT 2147.810 2994.620 2148.130 2994.680 ;
        RECT 2147.615 2994.480 2148.130 2994.620 ;
        RECT 2147.810 2994.420 2148.130 2994.480 ;
        RECT 2147.825 2946.680 2148.115 2946.725 ;
        RECT 2148.270 2946.680 2148.590 2946.740 ;
        RECT 2147.825 2946.540 2148.590 2946.680 ;
        RECT 2147.825 2946.495 2148.115 2946.540 ;
        RECT 2148.270 2946.480 2148.590 2946.540 ;
        RECT 2148.270 2912.340 2148.590 2912.400 ;
        RECT 2147.900 2912.200 2148.590 2912.340 ;
        RECT 2147.900 2911.720 2148.040 2912.200 ;
        RECT 2148.270 2912.140 2148.590 2912.200 ;
        RECT 2147.810 2911.460 2148.130 2911.720 ;
        RECT 2146.430 2815.580 2146.750 2815.840 ;
        RECT 2146.520 2815.160 2146.660 2815.580 ;
        RECT 2146.430 2814.900 2146.750 2815.160 ;
        RECT 2146.430 2801.160 2146.750 2801.220 ;
        RECT 2146.235 2801.020 2146.750 2801.160 ;
        RECT 2146.430 2800.960 2146.750 2801.020 ;
        RECT 2146.445 2753.220 2146.735 2753.265 ;
        RECT 2147.350 2753.220 2147.670 2753.280 ;
        RECT 2146.445 2753.080 2147.670 2753.220 ;
        RECT 2146.445 2753.035 2146.735 2753.080 ;
        RECT 2147.350 2753.020 2147.670 2753.080 ;
        RECT 2146.430 2718.200 2146.750 2718.260 ;
        RECT 2147.350 2718.200 2147.670 2718.260 ;
        RECT 2146.430 2718.060 2147.670 2718.200 ;
        RECT 2146.430 2718.000 2146.750 2718.060 ;
        RECT 2147.350 2718.000 2147.670 2718.060 ;
        RECT 2146.430 2670.260 2146.750 2670.320 ;
        RECT 2147.350 2670.260 2147.670 2670.320 ;
        RECT 2146.430 2670.120 2147.670 2670.260 ;
        RECT 2146.430 2670.060 2146.750 2670.120 ;
        RECT 2147.350 2670.060 2147.670 2670.120 ;
        RECT 2147.350 2622.120 2147.670 2622.380 ;
        RECT 2147.440 2621.980 2147.580 2622.120 ;
        RECT 2147.810 2621.980 2148.130 2622.040 ;
        RECT 2147.440 2621.840 2148.130 2621.980 ;
        RECT 2147.810 2621.780 2148.130 2621.840 ;
        RECT 2146.890 2560.100 2147.210 2560.160 ;
        RECT 2148.270 2560.100 2148.590 2560.160 ;
        RECT 2146.890 2559.960 2148.590 2560.100 ;
        RECT 2146.890 2559.900 2147.210 2559.960 ;
        RECT 2148.270 2559.900 2148.590 2559.960 ;
        RECT 2147.350 2511.820 2147.670 2511.880 ;
        RECT 2148.270 2511.820 2148.590 2511.880 ;
        RECT 2147.350 2511.680 2148.590 2511.820 ;
        RECT 2147.350 2511.620 2147.670 2511.680 ;
        RECT 2148.270 2511.620 2148.590 2511.680 ;
        RECT 2146.890 2463.200 2147.210 2463.260 ;
        RECT 2146.695 2463.060 2147.210 2463.200 ;
        RECT 2146.890 2463.000 2147.210 2463.060 ;
        RECT 2146.890 2428.860 2147.210 2428.920 ;
        RECT 2146.695 2428.720 2147.210 2428.860 ;
        RECT 2146.890 2428.660 2147.210 2428.720 ;
        RECT 2146.430 2380.580 2146.750 2380.640 ;
        RECT 2147.350 2380.580 2147.670 2380.640 ;
        RECT 2146.430 2380.440 2147.670 2380.580 ;
        RECT 2146.430 2380.380 2146.750 2380.440 ;
        RECT 2147.350 2380.380 2147.670 2380.440 ;
        RECT 2146.890 2366.640 2147.210 2366.700 ;
        RECT 2146.695 2366.500 2147.210 2366.640 ;
        RECT 2146.890 2366.440 2147.210 2366.500 ;
        RECT 2146.890 2331.960 2147.210 2332.020 ;
        RECT 2146.695 2331.820 2147.210 2331.960 ;
        RECT 2146.890 2331.760 2147.210 2331.820 ;
        RECT 2145.970 2235.540 2146.290 2235.800 ;
        RECT 2146.060 2235.400 2146.200 2235.540 ;
        RECT 2146.430 2235.400 2146.750 2235.460 ;
        RECT 2146.060 2235.260 2146.750 2235.400 ;
        RECT 2146.430 2235.200 2146.750 2235.260 ;
        RECT 2145.050 2221.800 2145.370 2221.860 ;
        RECT 2146.430 2221.800 2146.750 2221.860 ;
        RECT 2145.050 2221.660 2146.750 2221.800 ;
        RECT 2145.050 2221.600 2145.370 2221.660 ;
        RECT 2146.430 2221.600 2146.750 2221.660 ;
        RECT 2145.970 2138.980 2146.290 2139.240 ;
        RECT 2146.060 2138.840 2146.200 2138.980 ;
        RECT 2146.430 2138.840 2146.750 2138.900 ;
        RECT 2146.060 2138.700 2146.750 2138.840 ;
        RECT 2146.430 2138.640 2146.750 2138.700 ;
        RECT 2145.050 2125.240 2145.370 2125.300 ;
        RECT 2146.430 2125.240 2146.750 2125.300 ;
        RECT 2145.050 2125.100 2146.750 2125.240 ;
        RECT 2145.050 2125.040 2145.370 2125.100 ;
        RECT 2146.430 2125.040 2146.750 2125.100 ;
        RECT 2145.970 2042.420 2146.290 2042.680 ;
        RECT 2146.060 2041.940 2146.200 2042.420 ;
        RECT 2146.430 2041.940 2146.750 2042.000 ;
        RECT 2146.060 2041.800 2146.750 2041.940 ;
        RECT 2146.430 2041.740 2146.750 2041.800 ;
        RECT 2146.430 2028.340 2146.750 2028.400 ;
        RECT 2146.235 2028.200 2146.750 2028.340 ;
        RECT 2146.430 2028.140 2146.750 2028.200 ;
        RECT 2146.430 1994.000 2146.750 1994.060 ;
        RECT 2146.235 1993.860 2146.750 1994.000 ;
        RECT 2146.430 1993.800 2146.750 1993.860 ;
        RECT 2146.430 1945.860 2146.750 1946.120 ;
        RECT 2146.520 1945.440 2146.660 1945.860 ;
        RECT 2146.430 1945.180 2146.750 1945.440 ;
        RECT 2146.430 1897.440 2146.750 1897.500 ;
        RECT 2147.350 1897.440 2147.670 1897.500 ;
        RECT 2146.430 1897.300 2147.670 1897.440 ;
        RECT 2146.430 1897.240 2146.750 1897.300 ;
        RECT 2147.350 1897.240 2147.670 1897.300 ;
        RECT 2147.810 1787.620 2148.130 1787.680 ;
        RECT 2147.615 1787.480 2148.130 1787.620 ;
        RECT 2147.810 1787.420 2148.130 1787.480 ;
        RECT 2147.810 1766.880 2148.130 1766.940 ;
        RECT 2147.615 1766.740 2148.130 1766.880 ;
        RECT 2147.810 1766.680 2148.130 1766.740 ;
        RECT 2148.270 1766.200 2148.590 1766.260 ;
        RECT 2148.075 1766.060 2148.590 1766.200 ;
        RECT 2148.270 1766.000 2148.590 1766.060 ;
        RECT 2148.270 1703.980 2148.590 1704.040 ;
        RECT 2148.075 1703.840 2148.590 1703.980 ;
        RECT 2148.270 1703.780 2148.590 1703.840 ;
        RECT 2147.350 1628.500 2147.670 1628.560 ;
        RECT 2147.810 1628.500 2148.130 1628.560 ;
        RECT 2147.350 1628.360 2148.130 1628.500 ;
        RECT 2147.350 1628.300 2147.670 1628.360 ;
        RECT 2147.810 1628.300 2148.130 1628.360 ;
        RECT 2146.890 1594.160 2147.210 1594.220 ;
        RECT 2147.350 1594.160 2147.670 1594.220 ;
        RECT 2146.890 1594.020 2147.670 1594.160 ;
        RECT 2146.890 1593.960 2147.210 1594.020 ;
        RECT 2147.350 1593.960 2147.670 1594.020 ;
        RECT 2146.890 1559.820 2147.210 1559.880 ;
        RECT 2147.350 1559.820 2147.670 1559.880 ;
        RECT 2146.890 1559.680 2147.670 1559.820 ;
        RECT 2146.890 1559.620 2147.210 1559.680 ;
        RECT 2147.350 1559.620 2147.670 1559.680 ;
        RECT 2146.430 1511.200 2146.750 1511.260 ;
        RECT 2147.350 1511.200 2147.670 1511.260 ;
        RECT 2146.430 1511.060 2147.670 1511.200 ;
        RECT 2146.430 1511.000 2146.750 1511.060 ;
        RECT 2147.350 1511.000 2147.670 1511.060 ;
        RECT 2147.350 1448.980 2147.670 1449.040 ;
        RECT 2147.155 1448.840 2147.670 1448.980 ;
        RECT 2147.350 1448.780 2147.670 1448.840 ;
        RECT 2147.365 1401.040 2147.655 1401.085 ;
        RECT 2147.810 1401.040 2148.130 1401.100 ;
        RECT 2147.365 1400.900 2148.130 1401.040 ;
        RECT 2147.365 1400.855 2147.655 1400.900 ;
        RECT 2147.810 1400.840 2148.130 1400.900 ;
        RECT 2146.890 1374.520 2147.210 1374.580 ;
        RECT 2147.810 1374.520 2148.130 1374.580 ;
        RECT 2146.890 1374.380 2148.130 1374.520 ;
        RECT 2146.890 1374.320 2147.210 1374.380 ;
        RECT 2147.810 1374.320 2148.130 1374.380 ;
        RECT 2146.890 1352.420 2147.210 1352.480 ;
        RECT 2146.695 1352.280 2147.210 1352.420 ;
        RECT 2146.890 1352.220 2147.210 1352.280 ;
        RECT 2146.890 1317.740 2147.210 1317.800 ;
        RECT 2146.695 1317.600 2147.210 1317.740 ;
        RECT 2146.890 1317.540 2147.210 1317.600 ;
        RECT 2146.890 1304.140 2147.210 1304.200 ;
        RECT 2147.825 1304.140 2148.115 1304.185 ;
        RECT 2146.890 1304.000 2148.115 1304.140 ;
        RECT 2146.890 1303.940 2147.210 1304.000 ;
        RECT 2147.825 1303.955 2148.115 1304.000 ;
        RECT 2147.810 1269.800 2148.130 1269.860 ;
        RECT 2147.615 1269.660 2148.130 1269.800 ;
        RECT 2147.810 1269.600 2148.130 1269.660 ;
        RECT 2146.430 1173.380 2146.750 1173.640 ;
        RECT 2146.520 1172.960 2146.660 1173.380 ;
        RECT 2146.430 1172.700 2146.750 1172.960 ;
        RECT 2146.430 1158.960 2146.750 1159.020 ;
        RECT 2146.235 1158.820 2146.750 1158.960 ;
        RECT 2146.430 1158.760 2146.750 1158.820 ;
        RECT 2146.445 1111.020 2146.735 1111.065 ;
        RECT 2147.350 1111.020 2147.670 1111.080 ;
        RECT 2146.445 1110.880 2147.670 1111.020 ;
        RECT 2146.445 1110.835 2146.735 1110.880 ;
        RECT 2147.350 1110.820 2147.670 1110.880 ;
        RECT 2146.430 1076.000 2146.750 1076.060 ;
        RECT 2147.350 1076.000 2147.670 1076.060 ;
        RECT 2146.430 1075.860 2147.670 1076.000 ;
        RECT 2146.430 1075.800 2146.750 1075.860 ;
        RECT 2147.350 1075.800 2147.670 1075.860 ;
        RECT 2146.430 1028.060 2146.750 1028.120 ;
        RECT 2147.350 1028.060 2147.670 1028.120 ;
        RECT 2146.430 1027.920 2147.670 1028.060 ;
        RECT 2146.430 1027.860 2146.750 1027.920 ;
        RECT 2147.350 1027.860 2147.670 1027.920 ;
        RECT 2147.350 1014.120 2147.670 1014.180 ;
        RECT 2147.155 1013.980 2147.670 1014.120 ;
        RECT 2147.350 1013.920 2147.670 1013.980 ;
        RECT 2147.365 966.520 2147.655 966.565 ;
        RECT 2147.810 966.520 2148.130 966.580 ;
        RECT 2147.365 966.380 2148.130 966.520 ;
        RECT 2147.365 966.335 2147.655 966.380 ;
        RECT 2147.810 966.320 2148.130 966.380 ;
        RECT 2147.350 917.560 2147.670 917.620 ;
        RECT 2147.155 917.420 2147.670 917.560 ;
        RECT 2147.350 917.360 2147.670 917.420 ;
        RECT 2147.365 869.960 2147.655 870.005 ;
        RECT 2147.810 869.960 2148.130 870.020 ;
        RECT 2147.365 869.820 2148.130 869.960 ;
        RECT 2147.365 869.775 2147.655 869.820 ;
        RECT 2147.810 869.760 2148.130 869.820 ;
        RECT 2146.890 821.000 2147.210 821.060 ;
        RECT 2146.695 820.860 2147.210 821.000 ;
        RECT 2146.890 820.800 2147.210 820.860 ;
        RECT 2146.890 786.660 2147.210 786.720 ;
        RECT 2146.695 786.520 2147.210 786.660 ;
        RECT 2146.890 786.460 2147.210 786.520 ;
        RECT 2146.430 738.380 2146.750 738.440 ;
        RECT 2147.350 738.380 2147.670 738.440 ;
        RECT 2146.430 738.240 2147.670 738.380 ;
        RECT 2146.430 738.180 2146.750 738.240 ;
        RECT 2147.350 738.180 2147.670 738.240 ;
        RECT 2146.890 724.440 2147.210 724.500 ;
        RECT 2146.695 724.300 2147.210 724.440 ;
        RECT 2146.890 724.240 2147.210 724.300 ;
        RECT 2146.890 689.760 2147.210 689.820 ;
        RECT 2146.695 689.620 2147.210 689.760 ;
        RECT 2146.890 689.560 2147.210 689.620 ;
        RECT 2146.430 641.820 2146.750 641.880 ;
        RECT 2147.350 641.820 2147.670 641.880 ;
        RECT 2146.430 641.680 2147.670 641.820 ;
        RECT 2146.430 641.620 2146.750 641.680 ;
        RECT 2147.350 641.620 2147.670 641.680 ;
        RECT 2146.430 627.880 2146.750 627.940 ;
        RECT 2146.235 627.740 2146.750 627.880 ;
        RECT 2146.430 627.680 2146.750 627.740 ;
        RECT 2146.430 579.940 2146.750 580.000 ;
        RECT 2146.235 579.800 2146.750 579.940 ;
        RECT 2146.430 579.740 2146.750 579.800 ;
        RECT 2145.510 483.040 2145.830 483.100 ;
        RECT 2146.890 483.040 2147.210 483.100 ;
        RECT 2145.510 482.900 2147.210 483.040 ;
        RECT 2145.510 482.840 2145.830 482.900 ;
        RECT 2146.890 482.840 2147.210 482.900 ;
        RECT 2146.430 400.220 2146.750 400.480 ;
        RECT 2146.520 399.740 2146.660 400.220 ;
        RECT 2146.890 399.740 2147.210 399.800 ;
        RECT 2146.520 399.600 2147.210 399.740 ;
        RECT 2146.890 399.540 2147.210 399.600 ;
        RECT 2146.890 303.180 2147.210 303.240 ;
        RECT 2147.810 303.180 2148.130 303.240 ;
        RECT 2146.890 303.040 2148.130 303.180 ;
        RECT 2146.890 302.980 2147.210 303.040 ;
        RECT 2147.810 302.980 2148.130 303.040 ;
        RECT 1167.550 214.100 1167.870 214.160 ;
        RECT 2146.890 214.100 2147.210 214.160 ;
        RECT 1167.550 213.960 2147.210 214.100 ;
        RECT 1167.550 213.900 1167.870 213.960 ;
        RECT 2146.890 213.900 2147.210 213.960 ;
      LAYER via ;
        RECT 2146.920 3442.880 2147.180 3443.140 ;
        RECT 2149.220 3442.880 2149.480 3443.140 ;
        RECT 2146.460 3422.140 2146.720 3422.400 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.460 3056.640 2146.720 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 2146.920 3042.700 2147.180 3042.960 ;
        RECT 2147.840 3008.360 2148.100 3008.620 ;
        RECT 2147.840 2994.420 2148.100 2994.680 ;
        RECT 2148.300 2946.480 2148.560 2946.740 ;
        RECT 2148.300 2912.140 2148.560 2912.400 ;
        RECT 2147.840 2911.460 2148.100 2911.720 ;
        RECT 2146.460 2815.580 2146.720 2815.840 ;
        RECT 2146.460 2814.900 2146.720 2815.160 ;
        RECT 2146.460 2800.960 2146.720 2801.220 ;
        RECT 2147.380 2753.020 2147.640 2753.280 ;
        RECT 2146.460 2718.000 2146.720 2718.260 ;
        RECT 2147.380 2718.000 2147.640 2718.260 ;
        RECT 2146.460 2670.060 2146.720 2670.320 ;
        RECT 2147.380 2670.060 2147.640 2670.320 ;
        RECT 2147.380 2622.120 2147.640 2622.380 ;
        RECT 2147.840 2621.780 2148.100 2622.040 ;
        RECT 2146.920 2559.900 2147.180 2560.160 ;
        RECT 2148.300 2559.900 2148.560 2560.160 ;
        RECT 2147.380 2511.620 2147.640 2511.880 ;
        RECT 2148.300 2511.620 2148.560 2511.880 ;
        RECT 2146.920 2463.000 2147.180 2463.260 ;
        RECT 2146.920 2428.660 2147.180 2428.920 ;
        RECT 2146.460 2380.380 2146.720 2380.640 ;
        RECT 2147.380 2380.380 2147.640 2380.640 ;
        RECT 2146.920 2366.440 2147.180 2366.700 ;
        RECT 2146.920 2331.760 2147.180 2332.020 ;
        RECT 2146.000 2235.540 2146.260 2235.800 ;
        RECT 2146.460 2235.200 2146.720 2235.460 ;
        RECT 2145.080 2221.600 2145.340 2221.860 ;
        RECT 2146.460 2221.600 2146.720 2221.860 ;
        RECT 2146.000 2138.980 2146.260 2139.240 ;
        RECT 2146.460 2138.640 2146.720 2138.900 ;
        RECT 2145.080 2125.040 2145.340 2125.300 ;
        RECT 2146.460 2125.040 2146.720 2125.300 ;
        RECT 2146.000 2042.420 2146.260 2042.680 ;
        RECT 2146.460 2041.740 2146.720 2042.000 ;
        RECT 2146.460 2028.140 2146.720 2028.400 ;
        RECT 2146.460 1993.800 2146.720 1994.060 ;
        RECT 2146.460 1945.860 2146.720 1946.120 ;
        RECT 2146.460 1945.180 2146.720 1945.440 ;
        RECT 2146.460 1897.240 2146.720 1897.500 ;
        RECT 2147.380 1897.240 2147.640 1897.500 ;
        RECT 2147.840 1787.420 2148.100 1787.680 ;
        RECT 2147.840 1766.680 2148.100 1766.940 ;
        RECT 2148.300 1766.000 2148.560 1766.260 ;
        RECT 2148.300 1703.780 2148.560 1704.040 ;
        RECT 2147.380 1628.300 2147.640 1628.560 ;
        RECT 2147.840 1628.300 2148.100 1628.560 ;
        RECT 2146.920 1593.960 2147.180 1594.220 ;
        RECT 2147.380 1593.960 2147.640 1594.220 ;
        RECT 2146.920 1559.620 2147.180 1559.880 ;
        RECT 2147.380 1559.620 2147.640 1559.880 ;
        RECT 2146.460 1511.000 2146.720 1511.260 ;
        RECT 2147.380 1511.000 2147.640 1511.260 ;
        RECT 2147.380 1448.780 2147.640 1449.040 ;
        RECT 2147.840 1400.840 2148.100 1401.100 ;
        RECT 2146.920 1374.320 2147.180 1374.580 ;
        RECT 2147.840 1374.320 2148.100 1374.580 ;
        RECT 2146.920 1352.220 2147.180 1352.480 ;
        RECT 2146.920 1317.540 2147.180 1317.800 ;
        RECT 2146.920 1303.940 2147.180 1304.200 ;
        RECT 2147.840 1269.600 2148.100 1269.860 ;
        RECT 2146.460 1173.380 2146.720 1173.640 ;
        RECT 2146.460 1172.700 2146.720 1172.960 ;
        RECT 2146.460 1158.760 2146.720 1159.020 ;
        RECT 2147.380 1110.820 2147.640 1111.080 ;
        RECT 2146.460 1075.800 2146.720 1076.060 ;
        RECT 2147.380 1075.800 2147.640 1076.060 ;
        RECT 2146.460 1027.860 2146.720 1028.120 ;
        RECT 2147.380 1027.860 2147.640 1028.120 ;
        RECT 2147.380 1013.920 2147.640 1014.180 ;
        RECT 2147.840 966.320 2148.100 966.580 ;
        RECT 2147.380 917.360 2147.640 917.620 ;
        RECT 2147.840 869.760 2148.100 870.020 ;
        RECT 2146.920 820.800 2147.180 821.060 ;
        RECT 2146.920 786.460 2147.180 786.720 ;
        RECT 2146.460 738.180 2146.720 738.440 ;
        RECT 2147.380 738.180 2147.640 738.440 ;
        RECT 2146.920 724.240 2147.180 724.500 ;
        RECT 2146.920 689.560 2147.180 689.820 ;
        RECT 2146.460 641.620 2146.720 641.880 ;
        RECT 2147.380 641.620 2147.640 641.880 ;
        RECT 2146.460 627.680 2146.720 627.940 ;
        RECT 2146.460 579.740 2146.720 580.000 ;
        RECT 2145.540 482.840 2145.800 483.100 ;
        RECT 2146.920 482.840 2147.180 483.100 ;
        RECT 2146.460 400.220 2146.720 400.480 ;
        RECT 2146.920 399.540 2147.180 399.800 ;
        RECT 2146.920 302.980 2147.180 303.240 ;
        RECT 2147.840 302.980 2148.100 303.240 ;
        RECT 1167.580 213.900 1167.840 214.160 ;
        RECT 2146.920 213.900 2147.180 214.160 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3443.170 2149.420 3517.600 ;
        RECT 2146.920 3442.850 2147.180 3443.170 ;
        RECT 2149.220 3442.850 2149.480 3443.170 ;
        RECT 2146.980 3429.650 2147.120 3442.850 ;
        RECT 2146.520 3429.510 2147.120 3429.650 ;
        RECT 2146.520 3422.430 2146.660 3429.510 ;
        RECT 2146.460 3422.110 2146.720 3422.430 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3236.450 2147.580 3298.270 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3056.930 2147.580 3105.150 ;
        RECT 2146.460 3056.610 2146.720 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.520 3056.330 2146.660 3056.610 ;
        RECT 2146.520 3056.190 2147.120 3056.330 ;
        RECT 2146.980 3042.990 2147.120 3056.190 ;
        RECT 2146.920 3042.670 2147.180 3042.990 ;
        RECT 2147.840 3008.330 2148.100 3008.650 ;
        RECT 2147.900 2994.710 2148.040 3008.330 ;
        RECT 2147.840 2994.390 2148.100 2994.710 ;
        RECT 2148.300 2946.450 2148.560 2946.770 ;
        RECT 2148.360 2912.430 2148.500 2946.450 ;
        RECT 2148.300 2912.110 2148.560 2912.430 ;
        RECT 2147.840 2911.430 2148.100 2911.750 ;
        RECT 2147.900 2863.210 2148.040 2911.430 ;
        RECT 2146.980 2863.070 2148.040 2863.210 ;
        RECT 2146.980 2849.610 2147.120 2863.070 ;
        RECT 2146.520 2849.470 2147.120 2849.610 ;
        RECT 2146.520 2815.870 2146.660 2849.470 ;
        RECT 2146.460 2815.550 2146.720 2815.870 ;
        RECT 2146.460 2814.870 2146.720 2815.190 ;
        RECT 2146.520 2801.250 2146.660 2814.870 ;
        RECT 2146.460 2800.930 2146.720 2801.250 ;
        RECT 2147.380 2752.990 2147.640 2753.310 ;
        RECT 2147.440 2718.290 2147.580 2752.990 ;
        RECT 2146.460 2717.970 2146.720 2718.290 ;
        RECT 2147.380 2717.970 2147.640 2718.290 ;
        RECT 2146.520 2670.350 2146.660 2717.970 ;
        RECT 2146.460 2670.030 2146.720 2670.350 ;
        RECT 2147.380 2670.030 2147.640 2670.350 ;
        RECT 2147.440 2622.410 2147.580 2670.030 ;
        RECT 2147.380 2622.090 2147.640 2622.410 ;
        RECT 2147.840 2621.750 2148.100 2622.070 ;
        RECT 2147.900 2608.325 2148.040 2621.750 ;
        RECT 2146.910 2607.955 2147.190 2608.325 ;
        RECT 2147.830 2607.955 2148.110 2608.325 ;
        RECT 2146.980 2560.190 2147.120 2607.955 ;
        RECT 2146.920 2559.870 2147.180 2560.190 ;
        RECT 2148.300 2559.870 2148.560 2560.190 ;
        RECT 2148.360 2511.910 2148.500 2559.870 ;
        RECT 2147.380 2511.765 2147.640 2511.910 ;
        RECT 2145.990 2511.395 2146.270 2511.765 ;
        RECT 2147.370 2511.395 2147.650 2511.765 ;
        RECT 2148.300 2511.590 2148.560 2511.910 ;
        RECT 2146.060 2463.485 2146.200 2511.395 ;
        RECT 2145.990 2463.115 2146.270 2463.485 ;
        RECT 2146.910 2463.115 2147.190 2463.485 ;
        RECT 2146.920 2462.970 2147.180 2463.115 ;
        RECT 2146.920 2428.630 2147.180 2428.950 ;
        RECT 2146.980 2415.090 2147.120 2428.630 ;
        RECT 2146.980 2414.950 2147.580 2415.090 ;
        RECT 2147.440 2380.670 2147.580 2414.950 ;
        RECT 2146.460 2380.410 2146.720 2380.670 ;
        RECT 2146.460 2380.350 2147.120 2380.410 ;
        RECT 2147.380 2380.350 2147.640 2380.670 ;
        RECT 2146.520 2380.270 2147.120 2380.350 ;
        RECT 2146.980 2366.730 2147.120 2380.270 ;
        RECT 2146.920 2366.410 2147.180 2366.730 ;
        RECT 2146.920 2331.730 2147.180 2332.050 ;
        RECT 2146.980 2318.530 2147.120 2331.730 ;
        RECT 2146.980 2318.390 2147.580 2318.530 ;
        RECT 2147.440 2270.365 2147.580 2318.390 ;
        RECT 2145.990 2269.995 2146.270 2270.365 ;
        RECT 2147.370 2269.995 2147.650 2270.365 ;
        RECT 2146.060 2235.830 2146.200 2269.995 ;
        RECT 2146.000 2235.510 2146.260 2235.830 ;
        RECT 2146.460 2235.170 2146.720 2235.490 ;
        RECT 2146.520 2221.890 2146.660 2235.170 ;
        RECT 2145.080 2221.570 2145.340 2221.890 ;
        RECT 2146.460 2221.570 2146.720 2221.890 ;
        RECT 2145.140 2173.805 2145.280 2221.570 ;
        RECT 2145.070 2173.435 2145.350 2173.805 ;
        RECT 2145.990 2173.435 2146.270 2173.805 ;
        RECT 2146.060 2139.270 2146.200 2173.435 ;
        RECT 2146.000 2138.950 2146.260 2139.270 ;
        RECT 2146.460 2138.610 2146.720 2138.930 ;
        RECT 2146.520 2125.330 2146.660 2138.610 ;
        RECT 2145.080 2125.010 2145.340 2125.330 ;
        RECT 2146.460 2125.010 2146.720 2125.330 ;
        RECT 2145.140 2077.245 2145.280 2125.010 ;
        RECT 2145.070 2076.875 2145.350 2077.245 ;
        RECT 2145.990 2076.875 2146.270 2077.245 ;
        RECT 2146.060 2042.710 2146.200 2076.875 ;
        RECT 2146.000 2042.390 2146.260 2042.710 ;
        RECT 2146.460 2041.710 2146.720 2042.030 ;
        RECT 2146.520 2028.430 2146.660 2041.710 ;
        RECT 2146.460 2028.110 2146.720 2028.430 ;
        RECT 2146.460 1993.770 2146.720 1994.090 ;
        RECT 2146.520 1946.150 2146.660 1993.770 ;
        RECT 2146.460 1945.830 2146.720 1946.150 ;
        RECT 2146.460 1945.150 2146.720 1945.470 ;
        RECT 2146.520 1897.530 2146.660 1945.150 ;
        RECT 2146.460 1897.210 2146.720 1897.530 ;
        RECT 2147.380 1897.210 2147.640 1897.530 ;
        RECT 2147.440 1859.530 2147.580 1897.210 ;
        RECT 2147.440 1859.390 2148.040 1859.530 ;
        RECT 2147.900 1787.710 2148.040 1859.390 ;
        RECT 2147.840 1787.390 2148.100 1787.710 ;
        RECT 2147.840 1766.650 2148.100 1766.970 ;
        RECT 2147.900 1766.370 2148.040 1766.650 ;
        RECT 2147.900 1766.290 2148.500 1766.370 ;
        RECT 2147.900 1766.230 2148.560 1766.290 ;
        RECT 2148.300 1765.970 2148.560 1766.230 ;
        RECT 2148.300 1703.750 2148.560 1704.070 ;
        RECT 2148.360 1657.570 2148.500 1703.750 ;
        RECT 2147.900 1657.430 2148.500 1657.570 ;
        RECT 2147.900 1628.590 2148.040 1657.430 ;
        RECT 2147.380 1628.270 2147.640 1628.590 ;
        RECT 2147.840 1628.270 2148.100 1628.590 ;
        RECT 2147.440 1594.250 2147.580 1628.270 ;
        RECT 2146.920 1593.930 2147.180 1594.250 ;
        RECT 2147.380 1593.930 2147.640 1594.250 ;
        RECT 2146.980 1559.910 2147.120 1593.930 ;
        RECT 2146.920 1559.590 2147.180 1559.910 ;
        RECT 2147.380 1559.590 2147.640 1559.910 ;
        RECT 2147.440 1511.290 2147.580 1559.590 ;
        RECT 2146.460 1510.970 2146.720 1511.290 ;
        RECT 2147.380 1510.970 2147.640 1511.290 ;
        RECT 2146.520 1510.690 2146.660 1510.970 ;
        RECT 2146.520 1510.550 2147.120 1510.690 ;
        RECT 2146.980 1462.410 2147.120 1510.550 ;
        RECT 2146.980 1462.270 2147.580 1462.410 ;
        RECT 2147.440 1449.070 2147.580 1462.270 ;
        RECT 2147.380 1448.750 2147.640 1449.070 ;
        RECT 2147.840 1400.810 2148.100 1401.130 ;
        RECT 2147.900 1374.610 2148.040 1400.810 ;
        RECT 2146.920 1374.290 2147.180 1374.610 ;
        RECT 2147.840 1374.290 2148.100 1374.610 ;
        RECT 2146.980 1352.510 2147.120 1374.290 ;
        RECT 2146.920 1352.190 2147.180 1352.510 ;
        RECT 2146.920 1317.510 2147.180 1317.830 ;
        RECT 2146.980 1304.230 2147.120 1317.510 ;
        RECT 2146.920 1303.910 2147.180 1304.230 ;
        RECT 2147.840 1269.570 2148.100 1269.890 ;
        RECT 2147.900 1221.010 2148.040 1269.570 ;
        RECT 2146.980 1220.870 2148.040 1221.010 ;
        RECT 2146.980 1207.410 2147.120 1220.870 ;
        RECT 2146.520 1207.270 2147.120 1207.410 ;
        RECT 2146.520 1173.670 2146.660 1207.270 ;
        RECT 2146.460 1173.350 2146.720 1173.670 ;
        RECT 2146.460 1172.670 2146.720 1172.990 ;
        RECT 2146.520 1159.050 2146.660 1172.670 ;
        RECT 2146.460 1158.730 2146.720 1159.050 ;
        RECT 2147.380 1110.790 2147.640 1111.110 ;
        RECT 2147.440 1076.090 2147.580 1110.790 ;
        RECT 2146.460 1075.770 2146.720 1076.090 ;
        RECT 2147.380 1075.770 2147.640 1076.090 ;
        RECT 2146.520 1028.150 2146.660 1075.770 ;
        RECT 2146.460 1027.830 2146.720 1028.150 ;
        RECT 2147.380 1027.830 2147.640 1028.150 ;
        RECT 2147.440 1014.210 2147.580 1027.830 ;
        RECT 2147.380 1013.890 2147.640 1014.210 ;
        RECT 2147.840 966.290 2148.100 966.610 ;
        RECT 2147.900 931.330 2148.040 966.290 ;
        RECT 2147.440 931.190 2148.040 931.330 ;
        RECT 2147.440 917.650 2147.580 931.190 ;
        RECT 2147.380 917.330 2147.640 917.650 ;
        RECT 2147.840 869.730 2148.100 870.050 ;
        RECT 2147.900 834.770 2148.040 869.730 ;
        RECT 2146.980 834.630 2148.040 834.770 ;
        RECT 2146.980 821.090 2147.120 834.630 ;
        RECT 2146.920 820.770 2147.180 821.090 ;
        RECT 2146.920 786.430 2147.180 786.750 ;
        RECT 2146.980 772.890 2147.120 786.430 ;
        RECT 2146.980 772.750 2147.580 772.890 ;
        RECT 2147.440 738.470 2147.580 772.750 ;
        RECT 2146.460 738.210 2146.720 738.470 ;
        RECT 2146.460 738.150 2147.120 738.210 ;
        RECT 2147.380 738.150 2147.640 738.470 ;
        RECT 2146.520 738.070 2147.120 738.150 ;
        RECT 2146.980 724.530 2147.120 738.070 ;
        RECT 2146.920 724.210 2147.180 724.530 ;
        RECT 2146.920 689.530 2147.180 689.850 ;
        RECT 2146.980 676.330 2147.120 689.530 ;
        RECT 2146.980 676.190 2147.580 676.330 ;
        RECT 2147.440 641.910 2147.580 676.190 ;
        RECT 2146.460 641.590 2146.720 641.910 ;
        RECT 2147.380 641.590 2147.640 641.910 ;
        RECT 2146.520 627.970 2146.660 641.590 ;
        RECT 2146.460 627.650 2146.720 627.970 ;
        RECT 2146.460 579.710 2146.720 580.030 ;
        RECT 2146.520 545.090 2146.660 579.710 ;
        RECT 2146.520 544.950 2147.580 545.090 ;
        RECT 2147.440 507.010 2147.580 544.950 ;
        RECT 2146.980 506.870 2147.580 507.010 ;
        RECT 2146.980 483.130 2147.120 506.870 ;
        RECT 2145.540 482.810 2145.800 483.130 ;
        RECT 2146.920 482.810 2147.180 483.130 ;
        RECT 2145.600 435.045 2145.740 482.810 ;
        RECT 2145.530 434.675 2145.810 435.045 ;
        RECT 2146.450 434.675 2146.730 435.045 ;
        RECT 2146.520 400.510 2146.660 434.675 ;
        RECT 2146.460 400.190 2146.720 400.510 ;
        RECT 2146.920 399.510 2147.180 399.830 ;
        RECT 2146.980 352.650 2147.120 399.510 ;
        RECT 2146.980 352.510 2147.580 352.650 ;
        RECT 2147.440 351.290 2147.580 352.510 ;
        RECT 2146.520 351.150 2147.580 351.290 ;
        RECT 2146.520 337.805 2146.660 351.150 ;
        RECT 2146.450 337.435 2146.730 337.805 ;
        RECT 2147.830 337.435 2148.110 337.805 ;
        RECT 2147.900 303.270 2148.040 337.435 ;
        RECT 2146.920 302.950 2147.180 303.270 ;
        RECT 2147.840 302.950 2148.100 303.270 ;
        RECT 1167.530 216.000 1167.810 220.000 ;
        RECT 1167.640 214.190 1167.780 216.000 ;
        RECT 2146.980 214.190 2147.120 302.950 ;
        RECT 1167.580 213.870 1167.840 214.190 ;
        RECT 2146.920 213.870 2147.180 214.190 ;
      LAYER via2 ;
        RECT 2146.910 2608.000 2147.190 2608.280 ;
        RECT 2147.830 2608.000 2148.110 2608.280 ;
        RECT 2145.990 2511.440 2146.270 2511.720 ;
        RECT 2147.370 2511.440 2147.650 2511.720 ;
        RECT 2145.990 2463.160 2146.270 2463.440 ;
        RECT 2146.910 2463.160 2147.190 2463.440 ;
        RECT 2145.990 2270.040 2146.270 2270.320 ;
        RECT 2147.370 2270.040 2147.650 2270.320 ;
        RECT 2145.070 2173.480 2145.350 2173.760 ;
        RECT 2145.990 2173.480 2146.270 2173.760 ;
        RECT 2145.070 2076.920 2145.350 2077.200 ;
        RECT 2145.990 2076.920 2146.270 2077.200 ;
        RECT 2145.530 434.720 2145.810 435.000 ;
        RECT 2146.450 434.720 2146.730 435.000 ;
        RECT 2146.450 337.480 2146.730 337.760 ;
        RECT 2147.830 337.480 2148.110 337.760 ;
      LAYER met3 ;
        RECT 2146.885 2608.290 2147.215 2608.305 ;
        RECT 2147.805 2608.290 2148.135 2608.305 ;
        RECT 2146.885 2607.990 2148.135 2608.290 ;
        RECT 2146.885 2607.975 2147.215 2607.990 ;
        RECT 2147.805 2607.975 2148.135 2607.990 ;
        RECT 2145.965 2511.730 2146.295 2511.745 ;
        RECT 2147.345 2511.730 2147.675 2511.745 ;
        RECT 2145.965 2511.430 2147.675 2511.730 ;
        RECT 2145.965 2511.415 2146.295 2511.430 ;
        RECT 2147.345 2511.415 2147.675 2511.430 ;
        RECT 2145.965 2463.450 2146.295 2463.465 ;
        RECT 2146.885 2463.450 2147.215 2463.465 ;
        RECT 2145.965 2463.150 2147.215 2463.450 ;
        RECT 2145.965 2463.135 2146.295 2463.150 ;
        RECT 2146.885 2463.135 2147.215 2463.150 ;
        RECT 2145.965 2270.330 2146.295 2270.345 ;
        RECT 2147.345 2270.330 2147.675 2270.345 ;
        RECT 2145.965 2270.030 2147.675 2270.330 ;
        RECT 2145.965 2270.015 2146.295 2270.030 ;
        RECT 2147.345 2270.015 2147.675 2270.030 ;
        RECT 2145.045 2173.770 2145.375 2173.785 ;
        RECT 2145.965 2173.770 2146.295 2173.785 ;
        RECT 2145.045 2173.470 2146.295 2173.770 ;
        RECT 2145.045 2173.455 2145.375 2173.470 ;
        RECT 2145.965 2173.455 2146.295 2173.470 ;
        RECT 2145.045 2077.210 2145.375 2077.225 ;
        RECT 2145.965 2077.210 2146.295 2077.225 ;
        RECT 2145.045 2076.910 2146.295 2077.210 ;
        RECT 2145.045 2076.895 2145.375 2076.910 ;
        RECT 2145.965 2076.895 2146.295 2076.910 ;
        RECT 2145.505 435.010 2145.835 435.025 ;
        RECT 2146.425 435.010 2146.755 435.025 ;
        RECT 2145.505 434.710 2146.755 435.010 ;
        RECT 2145.505 434.695 2145.835 434.710 ;
        RECT 2146.425 434.695 2146.755 434.710 ;
        RECT 2146.425 337.770 2146.755 337.785 ;
        RECT 2147.805 337.770 2148.135 337.785 ;
        RECT 2146.425 337.470 2148.135 337.770 ;
        RECT 2146.425 337.455 2146.755 337.470 ;
        RECT 2147.805 337.455 2148.135 337.470 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1821.745 3332.765 1821.915 3380.875 ;
        RECT 1822.665 2753.065 1822.835 2767.175 ;
        RECT 1822.665 1787.465 1822.835 1801.235 ;
        RECT 1821.745 1690.565 1821.915 1738.675 ;
      LAYER mcon ;
        RECT 1821.745 3380.705 1821.915 3380.875 ;
        RECT 1822.665 2767.005 1822.835 2767.175 ;
        RECT 1822.665 1801.065 1822.835 1801.235 ;
        RECT 1821.745 1738.505 1821.915 1738.675 ;
      LAYER met1 ;
        RECT 1821.670 3380.860 1821.990 3380.920 ;
        RECT 1821.475 3380.720 1821.990 3380.860 ;
        RECT 1821.670 3380.660 1821.990 3380.720 ;
        RECT 1821.685 3332.920 1821.975 3332.965 ;
        RECT 1822.130 3332.920 1822.450 3332.980 ;
        RECT 1821.685 3332.780 1822.450 3332.920 ;
        RECT 1821.685 3332.735 1821.975 3332.780 ;
        RECT 1822.130 3332.720 1822.450 3332.780 ;
        RECT 1821.670 3270.700 1821.990 3270.760 ;
        RECT 1822.590 3270.700 1822.910 3270.760 ;
        RECT 1821.670 3270.560 1822.910 3270.700 ;
        RECT 1821.670 3270.500 1821.990 3270.560 ;
        RECT 1822.590 3270.500 1822.910 3270.560 ;
        RECT 1821.670 3174.140 1821.990 3174.200 ;
        RECT 1822.590 3174.140 1822.910 3174.200 ;
        RECT 1821.670 3174.000 1822.910 3174.140 ;
        RECT 1821.670 3173.940 1821.990 3174.000 ;
        RECT 1822.590 3173.940 1822.910 3174.000 ;
        RECT 1821.670 3077.580 1821.990 3077.640 ;
        RECT 1822.590 3077.580 1822.910 3077.640 ;
        RECT 1821.670 3077.440 1822.910 3077.580 ;
        RECT 1821.670 3077.380 1821.990 3077.440 ;
        RECT 1822.590 3077.380 1822.910 3077.440 ;
        RECT 1821.670 2981.020 1821.990 2981.080 ;
        RECT 1822.590 2981.020 1822.910 2981.080 ;
        RECT 1821.670 2980.880 1822.910 2981.020 ;
        RECT 1821.670 2980.820 1821.990 2980.880 ;
        RECT 1822.590 2980.820 1822.910 2980.880 ;
        RECT 1820.750 2946.340 1821.070 2946.400 ;
        RECT 1822.130 2946.340 1822.450 2946.400 ;
        RECT 1820.750 2946.200 1822.450 2946.340 ;
        RECT 1820.750 2946.140 1821.070 2946.200 ;
        RECT 1822.130 2946.140 1822.450 2946.200 ;
        RECT 1822.590 2767.160 1822.910 2767.220 ;
        RECT 1822.395 2767.020 1822.910 2767.160 ;
        RECT 1822.590 2766.960 1822.910 2767.020 ;
        RECT 1822.590 2753.220 1822.910 2753.280 ;
        RECT 1822.395 2753.080 1822.910 2753.220 ;
        RECT 1822.590 2753.020 1822.910 2753.080 ;
        RECT 1822.590 2719.020 1822.910 2719.280 ;
        RECT 1822.680 2718.880 1822.820 2719.020 ;
        RECT 1823.050 2718.880 1823.370 2718.940 ;
        RECT 1822.680 2718.740 1823.370 2718.880 ;
        RECT 1823.050 2718.680 1823.370 2718.740 ;
        RECT 1822.130 2656.660 1822.450 2656.720 ;
        RECT 1823.510 2656.660 1823.830 2656.720 ;
        RECT 1822.130 2656.520 1823.830 2656.660 ;
        RECT 1822.130 2656.460 1822.450 2656.520 ;
        RECT 1823.510 2656.460 1823.830 2656.520 ;
        RECT 1823.510 2622.660 1823.830 2622.720 ;
        RECT 1823.140 2622.520 1823.830 2622.660 ;
        RECT 1823.140 2622.040 1823.280 2622.520 ;
        RECT 1823.510 2622.460 1823.830 2622.520 ;
        RECT 1823.050 2621.780 1823.370 2622.040 ;
        RECT 1822.130 2560.100 1822.450 2560.160 ;
        RECT 1823.510 2560.100 1823.830 2560.160 ;
        RECT 1822.130 2559.960 1823.830 2560.100 ;
        RECT 1822.130 2559.900 1822.450 2559.960 ;
        RECT 1823.510 2559.900 1823.830 2559.960 ;
        RECT 1822.590 2511.820 1822.910 2511.880 ;
        RECT 1823.510 2511.820 1823.830 2511.880 ;
        RECT 1822.590 2511.680 1823.830 2511.820 ;
        RECT 1822.590 2511.620 1822.910 2511.680 ;
        RECT 1823.510 2511.620 1823.830 2511.680 ;
        RECT 1821.670 2401.320 1821.990 2401.380 ;
        RECT 1822.590 2401.320 1822.910 2401.380 ;
        RECT 1821.670 2401.180 1822.910 2401.320 ;
        RECT 1821.670 2401.120 1821.990 2401.180 ;
        RECT 1822.590 2401.120 1822.910 2401.180 ;
        RECT 1821.670 2304.760 1821.990 2304.820 ;
        RECT 1822.590 2304.760 1822.910 2304.820 ;
        RECT 1821.670 2304.620 1822.910 2304.760 ;
        RECT 1821.670 2304.560 1821.990 2304.620 ;
        RECT 1822.590 2304.560 1822.910 2304.620 ;
        RECT 1821.670 2208.200 1821.990 2208.260 ;
        RECT 1822.590 2208.200 1822.910 2208.260 ;
        RECT 1821.670 2208.060 1822.910 2208.200 ;
        RECT 1821.670 2208.000 1821.990 2208.060 ;
        RECT 1822.590 2208.000 1822.910 2208.060 ;
        RECT 1821.670 2111.640 1821.990 2111.700 ;
        RECT 1822.590 2111.640 1822.910 2111.700 ;
        RECT 1821.670 2111.500 1822.910 2111.640 ;
        RECT 1821.670 2111.440 1821.990 2111.500 ;
        RECT 1822.590 2111.440 1822.910 2111.500 ;
        RECT 1821.670 2015.080 1821.990 2015.140 ;
        RECT 1822.590 2015.080 1822.910 2015.140 ;
        RECT 1821.670 2014.940 1822.910 2015.080 ;
        RECT 1821.670 2014.880 1821.990 2014.940 ;
        RECT 1822.590 2014.880 1822.910 2014.940 ;
        RECT 1821.670 1918.520 1821.990 1918.580 ;
        RECT 1822.590 1918.520 1822.910 1918.580 ;
        RECT 1821.670 1918.380 1822.910 1918.520 ;
        RECT 1821.670 1918.320 1821.990 1918.380 ;
        RECT 1822.590 1918.320 1822.910 1918.380 ;
        RECT 1822.590 1801.220 1822.910 1801.280 ;
        RECT 1822.395 1801.080 1822.910 1801.220 ;
        RECT 1822.590 1801.020 1822.910 1801.080 ;
        RECT 1822.590 1787.620 1822.910 1787.680 ;
        RECT 1822.395 1787.480 1822.910 1787.620 ;
        RECT 1822.590 1787.420 1822.910 1787.480 ;
        RECT 1821.670 1738.660 1821.990 1738.720 ;
        RECT 1821.475 1738.520 1821.990 1738.660 ;
        RECT 1821.670 1738.460 1821.990 1738.520 ;
        RECT 1821.685 1690.720 1821.975 1690.765 ;
        RECT 1822.130 1690.720 1822.450 1690.780 ;
        RECT 1821.685 1690.580 1822.450 1690.720 ;
        RECT 1821.685 1690.535 1821.975 1690.580 ;
        RECT 1822.130 1690.520 1822.450 1690.580 ;
        RECT 1821.670 1628.500 1821.990 1628.560 ;
        RECT 1822.590 1628.500 1822.910 1628.560 ;
        RECT 1821.670 1628.360 1822.910 1628.500 ;
        RECT 1821.670 1628.300 1821.990 1628.360 ;
        RECT 1822.590 1628.300 1822.910 1628.360 ;
        RECT 1821.670 1531.940 1821.990 1532.000 ;
        RECT 1822.590 1531.940 1822.910 1532.000 ;
        RECT 1821.670 1531.800 1822.910 1531.940 ;
        RECT 1821.670 1531.740 1821.990 1531.800 ;
        RECT 1822.590 1531.740 1822.910 1531.800 ;
        RECT 1821.670 1435.380 1821.990 1435.440 ;
        RECT 1822.590 1435.380 1822.910 1435.440 ;
        RECT 1821.670 1435.240 1822.910 1435.380 ;
        RECT 1821.670 1435.180 1821.990 1435.240 ;
        RECT 1822.590 1435.180 1822.910 1435.240 ;
      LAYER via ;
        RECT 1821.700 3380.660 1821.960 3380.920 ;
        RECT 1822.160 3332.720 1822.420 3332.980 ;
        RECT 1821.700 3270.500 1821.960 3270.760 ;
        RECT 1822.620 3270.500 1822.880 3270.760 ;
        RECT 1821.700 3173.940 1821.960 3174.200 ;
        RECT 1822.620 3173.940 1822.880 3174.200 ;
        RECT 1821.700 3077.380 1821.960 3077.640 ;
        RECT 1822.620 3077.380 1822.880 3077.640 ;
        RECT 1821.700 2980.820 1821.960 2981.080 ;
        RECT 1822.620 2980.820 1822.880 2981.080 ;
        RECT 1820.780 2946.140 1821.040 2946.400 ;
        RECT 1822.160 2946.140 1822.420 2946.400 ;
        RECT 1822.620 2766.960 1822.880 2767.220 ;
        RECT 1822.620 2753.020 1822.880 2753.280 ;
        RECT 1822.620 2719.020 1822.880 2719.280 ;
        RECT 1823.080 2718.680 1823.340 2718.940 ;
        RECT 1822.160 2656.460 1822.420 2656.720 ;
        RECT 1823.540 2656.460 1823.800 2656.720 ;
        RECT 1823.540 2622.460 1823.800 2622.720 ;
        RECT 1823.080 2621.780 1823.340 2622.040 ;
        RECT 1822.160 2559.900 1822.420 2560.160 ;
        RECT 1823.540 2559.900 1823.800 2560.160 ;
        RECT 1822.620 2511.620 1822.880 2511.880 ;
        RECT 1823.540 2511.620 1823.800 2511.880 ;
        RECT 1821.700 2401.120 1821.960 2401.380 ;
        RECT 1822.620 2401.120 1822.880 2401.380 ;
        RECT 1821.700 2304.560 1821.960 2304.820 ;
        RECT 1822.620 2304.560 1822.880 2304.820 ;
        RECT 1821.700 2208.000 1821.960 2208.260 ;
        RECT 1822.620 2208.000 1822.880 2208.260 ;
        RECT 1821.700 2111.440 1821.960 2111.700 ;
        RECT 1822.620 2111.440 1822.880 2111.700 ;
        RECT 1821.700 2014.880 1821.960 2015.140 ;
        RECT 1822.620 2014.880 1822.880 2015.140 ;
        RECT 1821.700 1918.320 1821.960 1918.580 ;
        RECT 1822.620 1918.320 1822.880 1918.580 ;
        RECT 1822.620 1801.020 1822.880 1801.280 ;
        RECT 1822.620 1787.420 1822.880 1787.680 ;
        RECT 1821.700 1738.460 1821.960 1738.720 ;
        RECT 1822.160 1690.520 1822.420 1690.780 ;
        RECT 1821.700 1628.300 1821.960 1628.560 ;
        RECT 1822.620 1628.300 1822.880 1628.560 ;
        RECT 1821.700 1531.740 1821.960 1532.000 ;
        RECT 1822.620 1531.740 1822.880 1532.000 ;
        RECT 1821.700 1435.180 1821.960 1435.440 ;
        RECT 1822.620 1435.180 1822.880 1435.440 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3430.445 1825.580 3517.230 ;
        RECT 1825.370 3430.075 1825.650 3430.445 ;
        RECT 1822.610 3429.395 1822.890 3429.765 ;
        RECT 1822.680 3394.970 1822.820 3429.395 ;
        RECT 1821.760 3394.830 1822.820 3394.970 ;
        RECT 1821.760 3380.950 1821.900 3394.830 ;
        RECT 1821.700 3380.630 1821.960 3380.950 ;
        RECT 1822.160 3332.690 1822.420 3333.010 ;
        RECT 1822.220 3298.410 1822.360 3332.690 ;
        RECT 1822.220 3298.270 1822.820 3298.410 ;
        RECT 1822.680 3270.790 1822.820 3298.270 ;
        RECT 1821.700 3270.470 1821.960 3270.790 ;
        RECT 1822.620 3270.470 1822.880 3270.790 ;
        RECT 1821.760 3222.250 1821.900 3270.470 ;
        RECT 1821.760 3222.110 1822.820 3222.250 ;
        RECT 1822.680 3174.230 1822.820 3222.110 ;
        RECT 1821.700 3173.910 1821.960 3174.230 ;
        RECT 1822.620 3173.910 1822.880 3174.230 ;
        RECT 1821.760 3125.690 1821.900 3173.910 ;
        RECT 1821.760 3125.550 1822.820 3125.690 ;
        RECT 1822.680 3077.670 1822.820 3125.550 ;
        RECT 1821.700 3077.350 1821.960 3077.670 ;
        RECT 1822.620 3077.350 1822.880 3077.670 ;
        RECT 1821.760 3029.130 1821.900 3077.350 ;
        RECT 1821.760 3028.990 1822.820 3029.130 ;
        RECT 1822.680 2981.110 1822.820 3028.990 ;
        RECT 1821.700 2980.850 1821.960 2981.110 ;
        RECT 1821.700 2980.790 1822.360 2980.850 ;
        RECT 1822.620 2980.790 1822.880 2981.110 ;
        RECT 1821.760 2980.710 1822.360 2980.790 ;
        RECT 1822.220 2980.170 1822.360 2980.710 ;
        RECT 1822.220 2980.030 1822.820 2980.170 ;
        RECT 1822.680 2959.770 1822.820 2980.030 ;
        RECT 1822.220 2959.630 1822.820 2959.770 ;
        RECT 1822.220 2946.430 1822.360 2959.630 ;
        RECT 1820.780 2946.110 1821.040 2946.430 ;
        RECT 1822.160 2946.110 1822.420 2946.430 ;
        RECT 1820.840 2898.685 1820.980 2946.110 ;
        RECT 1820.770 2898.315 1821.050 2898.685 ;
        RECT 1821.690 2898.315 1821.970 2898.685 ;
        RECT 1821.760 2863.210 1821.900 2898.315 ;
        RECT 1821.760 2863.070 1822.360 2863.210 ;
        RECT 1822.220 2815.610 1822.360 2863.070 ;
        RECT 1822.220 2815.470 1822.820 2815.610 ;
        RECT 1822.680 2767.250 1822.820 2815.470 ;
        RECT 1822.620 2766.930 1822.880 2767.250 ;
        RECT 1822.620 2752.990 1822.880 2753.310 ;
        RECT 1822.680 2719.310 1822.820 2752.990 ;
        RECT 1822.620 2718.990 1822.880 2719.310 ;
        RECT 1823.080 2718.650 1823.340 2718.970 ;
        RECT 1823.140 2704.885 1823.280 2718.650 ;
        RECT 1822.150 2704.515 1822.430 2704.885 ;
        RECT 1823.070 2704.515 1823.350 2704.885 ;
        RECT 1822.220 2656.750 1822.360 2704.515 ;
        RECT 1822.160 2656.430 1822.420 2656.750 ;
        RECT 1823.540 2656.430 1823.800 2656.750 ;
        RECT 1823.600 2622.750 1823.740 2656.430 ;
        RECT 1823.540 2622.430 1823.800 2622.750 ;
        RECT 1823.080 2621.750 1823.340 2622.070 ;
        RECT 1823.140 2608.325 1823.280 2621.750 ;
        RECT 1822.150 2607.955 1822.430 2608.325 ;
        RECT 1823.070 2607.955 1823.350 2608.325 ;
        RECT 1822.220 2560.190 1822.360 2607.955 ;
        RECT 1822.160 2559.870 1822.420 2560.190 ;
        RECT 1823.540 2559.870 1823.800 2560.190 ;
        RECT 1823.600 2511.910 1823.740 2559.870 ;
        RECT 1822.620 2511.765 1822.880 2511.910 ;
        RECT 1821.230 2511.395 1821.510 2511.765 ;
        RECT 1822.610 2511.395 1822.890 2511.765 ;
        RECT 1823.540 2511.590 1823.800 2511.910 ;
        RECT 1821.300 2463.485 1821.440 2511.395 ;
        RECT 1821.230 2463.115 1821.510 2463.485 ;
        RECT 1822.150 2463.115 1822.430 2463.485 ;
        RECT 1822.220 2449.770 1822.360 2463.115 ;
        RECT 1822.220 2449.630 1822.820 2449.770 ;
        RECT 1822.680 2401.410 1822.820 2449.630 ;
        RECT 1821.700 2401.090 1821.960 2401.410 ;
        RECT 1822.620 2401.090 1822.880 2401.410 ;
        RECT 1821.760 2400.810 1821.900 2401.090 ;
        RECT 1821.760 2400.670 1822.360 2400.810 ;
        RECT 1822.220 2353.210 1822.360 2400.670 ;
        RECT 1822.220 2353.070 1822.820 2353.210 ;
        RECT 1822.680 2304.850 1822.820 2353.070 ;
        RECT 1821.700 2304.530 1821.960 2304.850 ;
        RECT 1822.620 2304.530 1822.880 2304.850 ;
        RECT 1821.760 2304.250 1821.900 2304.530 ;
        RECT 1821.760 2304.110 1822.360 2304.250 ;
        RECT 1822.220 2256.650 1822.360 2304.110 ;
        RECT 1822.220 2256.510 1822.820 2256.650 ;
        RECT 1822.680 2208.290 1822.820 2256.510 ;
        RECT 1821.700 2207.970 1821.960 2208.290 ;
        RECT 1822.620 2207.970 1822.880 2208.290 ;
        RECT 1821.760 2207.690 1821.900 2207.970 ;
        RECT 1821.760 2207.550 1822.360 2207.690 ;
        RECT 1822.220 2160.090 1822.360 2207.550 ;
        RECT 1822.220 2159.950 1822.820 2160.090 ;
        RECT 1822.680 2111.730 1822.820 2159.950 ;
        RECT 1821.700 2111.410 1821.960 2111.730 ;
        RECT 1822.620 2111.410 1822.880 2111.730 ;
        RECT 1821.760 2111.130 1821.900 2111.410 ;
        RECT 1821.760 2110.990 1822.360 2111.130 ;
        RECT 1822.220 2063.530 1822.360 2110.990 ;
        RECT 1822.220 2063.390 1822.820 2063.530 ;
        RECT 1822.680 2015.170 1822.820 2063.390 ;
        RECT 1821.700 2014.850 1821.960 2015.170 ;
        RECT 1822.620 2014.850 1822.880 2015.170 ;
        RECT 1821.760 2014.570 1821.900 2014.850 ;
        RECT 1821.760 2014.430 1822.360 2014.570 ;
        RECT 1822.220 1966.970 1822.360 2014.430 ;
        RECT 1822.220 1966.830 1822.820 1966.970 ;
        RECT 1822.680 1918.610 1822.820 1966.830 ;
        RECT 1821.700 1918.290 1821.960 1918.610 ;
        RECT 1822.620 1918.290 1822.880 1918.610 ;
        RECT 1821.760 1918.010 1821.900 1918.290 ;
        RECT 1821.760 1917.870 1822.360 1918.010 ;
        RECT 1822.220 1870.410 1822.360 1917.870 ;
        RECT 1822.220 1870.270 1822.820 1870.410 ;
        RECT 1822.680 1801.310 1822.820 1870.270 ;
        RECT 1822.620 1800.990 1822.880 1801.310 ;
        RECT 1822.620 1787.390 1822.880 1787.710 ;
        RECT 1822.680 1752.770 1822.820 1787.390 ;
        RECT 1821.760 1752.630 1822.820 1752.770 ;
        RECT 1821.760 1738.750 1821.900 1752.630 ;
        RECT 1821.700 1738.430 1821.960 1738.750 ;
        RECT 1822.160 1690.490 1822.420 1690.810 ;
        RECT 1822.220 1656.210 1822.360 1690.490 ;
        RECT 1822.220 1656.070 1822.820 1656.210 ;
        RECT 1822.680 1628.590 1822.820 1656.070 ;
        RECT 1821.700 1628.270 1821.960 1628.590 ;
        RECT 1822.620 1628.270 1822.880 1628.590 ;
        RECT 1821.760 1580.050 1821.900 1628.270 ;
        RECT 1821.760 1579.910 1822.820 1580.050 ;
        RECT 1822.680 1532.030 1822.820 1579.910 ;
        RECT 1821.700 1531.710 1821.960 1532.030 ;
        RECT 1822.620 1531.710 1822.880 1532.030 ;
        RECT 1821.760 1483.490 1821.900 1531.710 ;
        RECT 1821.760 1483.350 1822.820 1483.490 ;
        RECT 1822.680 1435.470 1822.820 1483.350 ;
        RECT 1821.700 1435.150 1821.960 1435.470 ;
        RECT 1822.620 1435.150 1822.880 1435.470 ;
        RECT 1821.760 1386.930 1821.900 1435.150 ;
        RECT 1821.760 1386.790 1822.820 1386.930 ;
        RECT 1822.680 1342.165 1822.820 1386.790 ;
        RECT 433.410 1341.795 433.690 1342.165 ;
        RECT 1822.610 1341.795 1822.890 1342.165 ;
        RECT 433.480 1325.025 433.620 1341.795 ;
        RECT 433.370 1321.025 433.650 1325.025 ;
      LAYER via2 ;
        RECT 1825.370 3430.120 1825.650 3430.400 ;
        RECT 1822.610 3429.440 1822.890 3429.720 ;
        RECT 1820.770 2898.360 1821.050 2898.640 ;
        RECT 1821.690 2898.360 1821.970 2898.640 ;
        RECT 1822.150 2704.560 1822.430 2704.840 ;
        RECT 1823.070 2704.560 1823.350 2704.840 ;
        RECT 1822.150 2608.000 1822.430 2608.280 ;
        RECT 1823.070 2608.000 1823.350 2608.280 ;
        RECT 1821.230 2511.440 1821.510 2511.720 ;
        RECT 1822.610 2511.440 1822.890 2511.720 ;
        RECT 1821.230 2463.160 1821.510 2463.440 ;
        RECT 1822.150 2463.160 1822.430 2463.440 ;
        RECT 433.410 1341.840 433.690 1342.120 ;
        RECT 1822.610 1341.840 1822.890 1342.120 ;
      LAYER met3 ;
        RECT 1825.345 3430.410 1825.675 3430.425 ;
        RECT 1821.910 3430.110 1825.675 3430.410 ;
        RECT 1821.910 3429.730 1822.210 3430.110 ;
        RECT 1825.345 3430.095 1825.675 3430.110 ;
        RECT 1822.585 3429.730 1822.915 3429.745 ;
        RECT 1821.910 3429.430 1822.915 3429.730 ;
        RECT 1822.585 3429.415 1822.915 3429.430 ;
        RECT 1820.745 2898.650 1821.075 2898.665 ;
        RECT 1821.665 2898.650 1821.995 2898.665 ;
        RECT 1820.745 2898.350 1821.995 2898.650 ;
        RECT 1820.745 2898.335 1821.075 2898.350 ;
        RECT 1821.665 2898.335 1821.995 2898.350 ;
        RECT 1822.125 2704.850 1822.455 2704.865 ;
        RECT 1823.045 2704.850 1823.375 2704.865 ;
        RECT 1822.125 2704.550 1823.375 2704.850 ;
        RECT 1822.125 2704.535 1822.455 2704.550 ;
        RECT 1823.045 2704.535 1823.375 2704.550 ;
        RECT 1822.125 2608.290 1822.455 2608.305 ;
        RECT 1823.045 2608.290 1823.375 2608.305 ;
        RECT 1822.125 2607.990 1823.375 2608.290 ;
        RECT 1822.125 2607.975 1822.455 2607.990 ;
        RECT 1823.045 2607.975 1823.375 2607.990 ;
        RECT 1821.205 2511.730 1821.535 2511.745 ;
        RECT 1822.585 2511.730 1822.915 2511.745 ;
        RECT 1821.205 2511.430 1822.915 2511.730 ;
        RECT 1821.205 2511.415 1821.535 2511.430 ;
        RECT 1822.585 2511.415 1822.915 2511.430 ;
        RECT 1821.205 2463.450 1821.535 2463.465 ;
        RECT 1822.125 2463.450 1822.455 2463.465 ;
        RECT 1821.205 2463.150 1822.455 2463.450 ;
        RECT 1821.205 2463.135 1821.535 2463.150 ;
        RECT 1822.125 2463.135 1822.455 2463.150 ;
        RECT 433.385 1342.130 433.715 1342.145 ;
        RECT 1822.585 1342.130 1822.915 1342.145 ;
        RECT 433.385 1341.830 1822.915 1342.130 ;
        RECT 433.385 1341.815 433.715 1341.830 ;
        RECT 1822.585 1341.815 1822.915 1341.830 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1499.285 3332.765 1499.455 3422.355 ;
        RECT 1498.365 3008.405 1498.535 3042.915 ;
        RECT 1499.285 2946.525 1499.455 2994.635 ;
        RECT 1498.365 2428.705 1498.535 2463.215 ;
        RECT 1498.365 2331.805 1498.535 2366.655 ;
        RECT 1497.445 2201.245 1497.615 2249.355 ;
        RECT 1497.445 2118.285 1497.615 2184.075 ;
        RECT 1497.905 1945.225 1498.075 1959.675 ;
        RECT 1499.285 1780.665 1499.455 1787.635 ;
        RECT 1499.285 1683.765 1499.455 1773.355 ;
        RECT 1498.365 1449.165 1498.535 1497.275 ;
        RECT 1498.365 966.365 1498.535 1014.135 ;
        RECT 1498.365 496.485 1498.535 507.195 ;
        RECT 1498.365 386.325 1498.535 434.775 ;
        RECT 1498.365 304.725 1498.535 337.875 ;
      LAYER mcon ;
        RECT 1499.285 3422.185 1499.455 3422.355 ;
        RECT 1498.365 3042.745 1498.535 3042.915 ;
        RECT 1499.285 2994.465 1499.455 2994.635 ;
        RECT 1498.365 2463.045 1498.535 2463.215 ;
        RECT 1498.365 2366.485 1498.535 2366.655 ;
        RECT 1497.445 2249.185 1497.615 2249.355 ;
        RECT 1497.445 2183.905 1497.615 2184.075 ;
        RECT 1497.905 1959.505 1498.075 1959.675 ;
        RECT 1499.285 1787.465 1499.455 1787.635 ;
        RECT 1499.285 1773.185 1499.455 1773.355 ;
        RECT 1498.365 1497.105 1498.535 1497.275 ;
        RECT 1498.365 1013.965 1498.535 1014.135 ;
        RECT 1498.365 507.025 1498.535 507.195 ;
        RECT 1498.365 434.605 1498.535 434.775 ;
        RECT 1498.365 337.705 1498.535 337.875 ;
      LAYER met1 ;
        RECT 1498.290 3443.080 1498.610 3443.140 ;
        RECT 1500.590 3443.080 1500.910 3443.140 ;
        RECT 1498.290 3442.940 1500.910 3443.080 ;
        RECT 1498.290 3442.880 1498.610 3442.940 ;
        RECT 1500.590 3442.880 1500.910 3442.940 ;
        RECT 1497.830 3422.340 1498.150 3422.400 ;
        RECT 1499.225 3422.340 1499.515 3422.385 ;
        RECT 1497.830 3422.200 1499.515 3422.340 ;
        RECT 1497.830 3422.140 1498.150 3422.200 ;
        RECT 1499.225 3422.155 1499.515 3422.200 ;
        RECT 1499.225 3332.920 1499.515 3332.965 ;
        RECT 1499.670 3332.920 1499.990 3332.980 ;
        RECT 1499.225 3332.780 1499.990 3332.920 ;
        RECT 1499.225 3332.735 1499.515 3332.780 ;
        RECT 1499.670 3332.720 1499.990 3332.780 ;
        RECT 1498.290 3236.360 1498.610 3236.420 ;
        RECT 1498.750 3236.360 1499.070 3236.420 ;
        RECT 1498.290 3236.220 1499.070 3236.360 ;
        RECT 1498.290 3236.160 1498.610 3236.220 ;
        RECT 1498.750 3236.160 1499.070 3236.220 ;
        RECT 1498.290 3202.020 1498.610 3202.080 ;
        RECT 1498.750 3202.020 1499.070 3202.080 ;
        RECT 1498.290 3201.880 1499.070 3202.020 ;
        RECT 1498.290 3201.820 1498.610 3201.880 ;
        RECT 1498.750 3201.820 1499.070 3201.880 ;
        RECT 1497.830 3153.400 1498.150 3153.460 ;
        RECT 1498.750 3153.400 1499.070 3153.460 ;
        RECT 1497.830 3153.260 1499.070 3153.400 ;
        RECT 1497.830 3153.200 1498.150 3153.260 ;
        RECT 1498.750 3153.200 1499.070 3153.260 ;
        RECT 1497.830 3056.840 1498.150 3056.900 ;
        RECT 1498.750 3056.840 1499.070 3056.900 ;
        RECT 1497.830 3056.700 1499.070 3056.840 ;
        RECT 1497.830 3056.640 1498.150 3056.700 ;
        RECT 1498.750 3056.640 1499.070 3056.700 ;
        RECT 1498.290 3042.900 1498.610 3042.960 ;
        RECT 1498.095 3042.760 1498.610 3042.900 ;
        RECT 1498.290 3042.700 1498.610 3042.760 ;
        RECT 1498.305 3008.560 1498.595 3008.605 ;
        RECT 1499.210 3008.560 1499.530 3008.620 ;
        RECT 1498.305 3008.420 1499.530 3008.560 ;
        RECT 1498.305 3008.375 1498.595 3008.420 ;
        RECT 1499.210 3008.360 1499.530 3008.420 ;
        RECT 1499.210 2994.620 1499.530 2994.680 ;
        RECT 1499.015 2994.480 1499.530 2994.620 ;
        RECT 1499.210 2994.420 1499.530 2994.480 ;
        RECT 1499.225 2946.680 1499.515 2946.725 ;
        RECT 1499.670 2946.680 1499.990 2946.740 ;
        RECT 1499.225 2946.540 1499.990 2946.680 ;
        RECT 1499.225 2946.495 1499.515 2946.540 ;
        RECT 1499.670 2946.480 1499.990 2946.540 ;
        RECT 1499.670 2912.340 1499.990 2912.400 ;
        RECT 1499.300 2912.200 1499.990 2912.340 ;
        RECT 1499.300 2911.720 1499.440 2912.200 ;
        RECT 1499.670 2912.140 1499.990 2912.200 ;
        RECT 1499.210 2911.460 1499.530 2911.720 ;
        RECT 1497.370 2753.220 1497.690 2753.280 ;
        RECT 1498.290 2753.220 1498.610 2753.280 ;
        RECT 1497.370 2753.080 1498.610 2753.220 ;
        RECT 1497.370 2753.020 1497.690 2753.080 ;
        RECT 1498.290 2753.020 1498.610 2753.080 ;
        RECT 1496.450 2718.540 1496.770 2718.600 ;
        RECT 1497.370 2718.540 1497.690 2718.600 ;
        RECT 1496.450 2718.400 1497.690 2718.540 ;
        RECT 1496.450 2718.340 1496.770 2718.400 ;
        RECT 1497.370 2718.340 1497.690 2718.400 ;
        RECT 1497.830 2656.660 1498.150 2656.720 ;
        RECT 1498.750 2656.660 1499.070 2656.720 ;
        RECT 1497.830 2656.520 1499.070 2656.660 ;
        RECT 1497.830 2656.460 1498.150 2656.520 ;
        RECT 1498.750 2656.460 1499.070 2656.520 ;
        RECT 1498.750 2622.120 1499.070 2622.380 ;
        RECT 1498.840 2621.980 1498.980 2622.120 ;
        RECT 1499.210 2621.980 1499.530 2622.040 ;
        RECT 1498.840 2621.840 1499.530 2621.980 ;
        RECT 1499.210 2621.780 1499.530 2621.840 ;
        RECT 1498.290 2560.100 1498.610 2560.160 ;
        RECT 1499.670 2560.100 1499.990 2560.160 ;
        RECT 1498.290 2559.960 1499.990 2560.100 ;
        RECT 1498.290 2559.900 1498.610 2559.960 ;
        RECT 1499.670 2559.900 1499.990 2559.960 ;
        RECT 1498.750 2511.820 1499.070 2511.880 ;
        RECT 1499.670 2511.820 1499.990 2511.880 ;
        RECT 1498.750 2511.680 1499.990 2511.820 ;
        RECT 1498.750 2511.620 1499.070 2511.680 ;
        RECT 1499.670 2511.620 1499.990 2511.680 ;
        RECT 1498.290 2463.200 1498.610 2463.260 ;
        RECT 1498.095 2463.060 1498.610 2463.200 ;
        RECT 1498.290 2463.000 1498.610 2463.060 ;
        RECT 1498.290 2428.860 1498.610 2428.920 ;
        RECT 1498.095 2428.720 1498.610 2428.860 ;
        RECT 1498.290 2428.660 1498.610 2428.720 ;
        RECT 1497.830 2380.580 1498.150 2380.640 ;
        RECT 1498.750 2380.580 1499.070 2380.640 ;
        RECT 1497.830 2380.440 1499.070 2380.580 ;
        RECT 1497.830 2380.380 1498.150 2380.440 ;
        RECT 1498.750 2380.380 1499.070 2380.440 ;
        RECT 1498.290 2366.640 1498.610 2366.700 ;
        RECT 1498.095 2366.500 1498.610 2366.640 ;
        RECT 1498.290 2366.440 1498.610 2366.500 ;
        RECT 1498.290 2331.960 1498.610 2332.020 ;
        RECT 1498.095 2331.820 1498.610 2331.960 ;
        RECT 1498.290 2331.760 1498.610 2331.820 ;
        RECT 1496.910 2304.420 1497.230 2304.480 ;
        RECT 1498.750 2304.420 1499.070 2304.480 ;
        RECT 1496.910 2304.280 1499.070 2304.420 ;
        RECT 1496.910 2304.220 1497.230 2304.280 ;
        RECT 1498.750 2304.220 1499.070 2304.280 ;
        RECT 1497.370 2249.340 1497.690 2249.400 ;
        RECT 1497.175 2249.200 1497.690 2249.340 ;
        RECT 1497.370 2249.140 1497.690 2249.200 ;
        RECT 1497.385 2201.400 1497.675 2201.445 ;
        RECT 1497.830 2201.400 1498.150 2201.460 ;
        RECT 1497.385 2201.260 1498.150 2201.400 ;
        RECT 1497.385 2201.215 1497.675 2201.260 ;
        RECT 1497.830 2201.200 1498.150 2201.260 ;
        RECT 1497.385 2184.060 1497.675 2184.105 ;
        RECT 1497.830 2184.060 1498.150 2184.120 ;
        RECT 1497.385 2183.920 1498.150 2184.060 ;
        RECT 1497.385 2183.875 1497.675 2183.920 ;
        RECT 1497.830 2183.860 1498.150 2183.920 ;
        RECT 1497.385 2118.440 1497.675 2118.485 ;
        RECT 1497.830 2118.440 1498.150 2118.500 ;
        RECT 1497.385 2118.300 1498.150 2118.440 ;
        RECT 1497.385 2118.255 1497.675 2118.300 ;
        RECT 1497.830 2118.240 1498.150 2118.300 ;
        RECT 1497.830 2111.300 1498.150 2111.360 ;
        RECT 1498.750 2111.300 1499.070 2111.360 ;
        RECT 1497.830 2111.160 1499.070 2111.300 ;
        RECT 1497.830 2111.100 1498.150 2111.160 ;
        RECT 1498.750 2111.100 1499.070 2111.160 ;
        RECT 1497.370 2063.020 1497.690 2063.080 ;
        RECT 1497.830 2063.020 1498.150 2063.080 ;
        RECT 1497.370 2062.880 1498.150 2063.020 ;
        RECT 1497.370 2062.820 1497.690 2062.880 ;
        RECT 1497.830 2062.820 1498.150 2062.880 ;
        RECT 1495.990 2007.940 1496.310 2008.000 ;
        RECT 1497.830 2007.940 1498.150 2008.000 ;
        RECT 1495.990 2007.800 1498.150 2007.940 ;
        RECT 1495.990 2007.740 1496.310 2007.800 ;
        RECT 1497.830 2007.740 1498.150 2007.800 ;
        RECT 1496.910 1959.660 1497.230 1959.720 ;
        RECT 1497.845 1959.660 1498.135 1959.705 ;
        RECT 1496.910 1959.520 1498.135 1959.660 ;
        RECT 1496.910 1959.460 1497.230 1959.520 ;
        RECT 1497.845 1959.475 1498.135 1959.520 ;
        RECT 1497.830 1945.380 1498.150 1945.440 ;
        RECT 1497.635 1945.240 1498.150 1945.380 ;
        RECT 1497.830 1945.180 1498.150 1945.240 ;
        RECT 1497.830 1897.440 1498.150 1897.500 ;
        RECT 1498.750 1897.440 1499.070 1897.500 ;
        RECT 1497.830 1897.300 1499.070 1897.440 ;
        RECT 1497.830 1897.240 1498.150 1897.300 ;
        RECT 1498.750 1897.240 1499.070 1897.300 ;
        RECT 1499.210 1787.620 1499.530 1787.680 ;
        RECT 1499.015 1787.480 1499.530 1787.620 ;
        RECT 1499.210 1787.420 1499.530 1787.480 ;
        RECT 1498.750 1780.820 1499.070 1780.880 ;
        RECT 1499.225 1780.820 1499.515 1780.865 ;
        RECT 1498.750 1780.680 1499.515 1780.820 ;
        RECT 1498.750 1780.620 1499.070 1780.680 ;
        RECT 1499.225 1780.635 1499.515 1780.680 ;
        RECT 1499.210 1773.340 1499.530 1773.400 ;
        RECT 1499.015 1773.200 1499.530 1773.340 ;
        RECT 1499.210 1773.140 1499.530 1773.200 ;
        RECT 1499.225 1683.920 1499.515 1683.965 ;
        RECT 1499.670 1683.920 1499.990 1683.980 ;
        RECT 1499.225 1683.780 1499.990 1683.920 ;
        RECT 1499.225 1683.735 1499.515 1683.780 ;
        RECT 1499.670 1683.720 1499.990 1683.780 ;
        RECT 1498.750 1635.640 1499.070 1635.700 ;
        RECT 1499.210 1635.640 1499.530 1635.700 ;
        RECT 1498.750 1635.500 1499.530 1635.640 ;
        RECT 1498.750 1635.440 1499.070 1635.500 ;
        RECT 1499.210 1635.440 1499.530 1635.500 ;
        RECT 1498.290 1594.160 1498.610 1594.220 ;
        RECT 1498.750 1594.160 1499.070 1594.220 ;
        RECT 1498.290 1594.020 1499.070 1594.160 ;
        RECT 1498.290 1593.960 1498.610 1594.020 ;
        RECT 1498.750 1593.960 1499.070 1594.020 ;
        RECT 1498.290 1559.820 1498.610 1559.880 ;
        RECT 1498.750 1559.820 1499.070 1559.880 ;
        RECT 1498.290 1559.680 1499.070 1559.820 ;
        RECT 1498.290 1559.620 1498.610 1559.680 ;
        RECT 1498.750 1559.620 1499.070 1559.680 ;
        RECT 1497.830 1511.200 1498.150 1511.260 ;
        RECT 1498.750 1511.200 1499.070 1511.260 ;
        RECT 1497.830 1511.060 1499.070 1511.200 ;
        RECT 1497.830 1511.000 1498.150 1511.060 ;
        RECT 1498.750 1511.000 1499.070 1511.060 ;
        RECT 1498.290 1497.260 1498.610 1497.320 ;
        RECT 1498.095 1497.120 1498.610 1497.260 ;
        RECT 1498.290 1497.060 1498.610 1497.120 ;
        RECT 1498.305 1449.320 1498.595 1449.365 ;
        RECT 1498.750 1449.320 1499.070 1449.380 ;
        RECT 1498.305 1449.180 1499.070 1449.320 ;
        RECT 1498.305 1449.135 1498.595 1449.180 ;
        RECT 1498.750 1449.120 1499.070 1449.180 ;
        RECT 1497.370 1304.140 1497.690 1304.200 ;
        RECT 1498.290 1304.140 1498.610 1304.200 ;
        RECT 1497.370 1304.000 1498.610 1304.140 ;
        RECT 1497.370 1303.940 1497.690 1304.000 ;
        RECT 1498.290 1303.940 1498.610 1304.000 ;
        RECT 1497.370 1159.300 1497.690 1159.360 ;
        RECT 1498.750 1159.300 1499.070 1159.360 ;
        RECT 1497.370 1159.160 1499.070 1159.300 ;
        RECT 1497.370 1159.100 1497.690 1159.160 ;
        RECT 1498.750 1159.100 1499.070 1159.160 ;
        RECT 1497.370 1063.080 1497.690 1063.140 ;
        RECT 1498.750 1063.080 1499.070 1063.140 ;
        RECT 1497.370 1062.940 1499.070 1063.080 ;
        RECT 1497.370 1062.880 1497.690 1062.940 ;
        RECT 1498.750 1062.880 1499.070 1062.940 ;
        RECT 1498.290 1014.120 1498.610 1014.180 ;
        RECT 1498.095 1013.980 1498.610 1014.120 ;
        RECT 1498.290 1013.920 1498.610 1013.980 ;
        RECT 1498.305 966.520 1498.595 966.565 ;
        RECT 1498.750 966.520 1499.070 966.580 ;
        RECT 1498.305 966.380 1499.070 966.520 ;
        RECT 1498.305 966.335 1498.595 966.380 ;
        RECT 1498.750 966.320 1499.070 966.380 ;
        RECT 1497.370 869.960 1497.690 870.020 ;
        RECT 1498.750 869.960 1499.070 870.020 ;
        RECT 1497.370 869.820 1499.070 869.960 ;
        RECT 1497.370 869.760 1497.690 869.820 ;
        RECT 1498.750 869.760 1499.070 869.820 ;
        RECT 1497.370 821.000 1497.690 821.060 ;
        RECT 1498.290 821.000 1498.610 821.060 ;
        RECT 1497.370 820.860 1498.610 821.000 ;
        RECT 1497.370 820.800 1497.690 820.860 ;
        RECT 1498.290 820.800 1498.610 820.860 ;
        RECT 1498.290 507.180 1498.610 507.240 ;
        RECT 1498.095 507.040 1498.610 507.180 ;
        RECT 1498.290 506.980 1498.610 507.040 ;
        RECT 1498.290 496.640 1498.610 496.700 ;
        RECT 1498.095 496.500 1498.610 496.640 ;
        RECT 1498.290 496.440 1498.610 496.500 ;
        RECT 1498.290 434.760 1498.610 434.820 ;
        RECT 1498.095 434.620 1498.610 434.760 ;
        RECT 1498.290 434.560 1498.610 434.620 ;
        RECT 1498.290 386.480 1498.610 386.540 ;
        RECT 1498.095 386.340 1498.610 386.480 ;
        RECT 1498.290 386.280 1498.610 386.340 ;
        RECT 1498.290 337.860 1498.610 337.920 ;
        RECT 1498.095 337.720 1498.610 337.860 ;
        RECT 1498.290 337.660 1498.610 337.720 ;
        RECT 1498.290 304.880 1498.610 304.940 ;
        RECT 1498.095 304.740 1498.610 304.880 ;
        RECT 1498.290 304.680 1498.610 304.740 ;
        RECT 406.710 199.480 407.030 199.540 ;
        RECT 1498.750 199.480 1499.070 199.540 ;
        RECT 406.710 199.340 1499.070 199.480 ;
        RECT 406.710 199.280 407.030 199.340 ;
        RECT 1498.750 199.280 1499.070 199.340 ;
      LAYER via ;
        RECT 1498.320 3442.880 1498.580 3443.140 ;
        RECT 1500.620 3442.880 1500.880 3443.140 ;
        RECT 1497.860 3422.140 1498.120 3422.400 ;
        RECT 1499.700 3332.720 1499.960 3332.980 ;
        RECT 1498.320 3236.160 1498.580 3236.420 ;
        RECT 1498.780 3236.160 1499.040 3236.420 ;
        RECT 1498.320 3201.820 1498.580 3202.080 ;
        RECT 1498.780 3201.820 1499.040 3202.080 ;
        RECT 1497.860 3153.200 1498.120 3153.460 ;
        RECT 1498.780 3153.200 1499.040 3153.460 ;
        RECT 1497.860 3056.640 1498.120 3056.900 ;
        RECT 1498.780 3056.640 1499.040 3056.900 ;
        RECT 1498.320 3042.700 1498.580 3042.960 ;
        RECT 1499.240 3008.360 1499.500 3008.620 ;
        RECT 1499.240 2994.420 1499.500 2994.680 ;
        RECT 1499.700 2946.480 1499.960 2946.740 ;
        RECT 1499.700 2912.140 1499.960 2912.400 ;
        RECT 1499.240 2911.460 1499.500 2911.720 ;
        RECT 1497.400 2753.020 1497.660 2753.280 ;
        RECT 1498.320 2753.020 1498.580 2753.280 ;
        RECT 1496.480 2718.340 1496.740 2718.600 ;
        RECT 1497.400 2718.340 1497.660 2718.600 ;
        RECT 1497.860 2656.460 1498.120 2656.720 ;
        RECT 1498.780 2656.460 1499.040 2656.720 ;
        RECT 1498.780 2622.120 1499.040 2622.380 ;
        RECT 1499.240 2621.780 1499.500 2622.040 ;
        RECT 1498.320 2559.900 1498.580 2560.160 ;
        RECT 1499.700 2559.900 1499.960 2560.160 ;
        RECT 1498.780 2511.620 1499.040 2511.880 ;
        RECT 1499.700 2511.620 1499.960 2511.880 ;
        RECT 1498.320 2463.000 1498.580 2463.260 ;
        RECT 1498.320 2428.660 1498.580 2428.920 ;
        RECT 1497.860 2380.380 1498.120 2380.640 ;
        RECT 1498.780 2380.380 1499.040 2380.640 ;
        RECT 1498.320 2366.440 1498.580 2366.700 ;
        RECT 1498.320 2331.760 1498.580 2332.020 ;
        RECT 1496.940 2304.220 1497.200 2304.480 ;
        RECT 1498.780 2304.220 1499.040 2304.480 ;
        RECT 1497.400 2249.140 1497.660 2249.400 ;
        RECT 1497.860 2201.200 1498.120 2201.460 ;
        RECT 1497.860 2183.860 1498.120 2184.120 ;
        RECT 1497.860 2118.240 1498.120 2118.500 ;
        RECT 1497.860 2111.100 1498.120 2111.360 ;
        RECT 1498.780 2111.100 1499.040 2111.360 ;
        RECT 1497.400 2062.820 1497.660 2063.080 ;
        RECT 1497.860 2062.820 1498.120 2063.080 ;
        RECT 1496.020 2007.740 1496.280 2008.000 ;
        RECT 1497.860 2007.740 1498.120 2008.000 ;
        RECT 1496.940 1959.460 1497.200 1959.720 ;
        RECT 1497.860 1945.180 1498.120 1945.440 ;
        RECT 1497.860 1897.240 1498.120 1897.500 ;
        RECT 1498.780 1897.240 1499.040 1897.500 ;
        RECT 1499.240 1787.420 1499.500 1787.680 ;
        RECT 1498.780 1780.620 1499.040 1780.880 ;
        RECT 1499.240 1773.140 1499.500 1773.400 ;
        RECT 1499.700 1683.720 1499.960 1683.980 ;
        RECT 1498.780 1635.440 1499.040 1635.700 ;
        RECT 1499.240 1635.440 1499.500 1635.700 ;
        RECT 1498.320 1593.960 1498.580 1594.220 ;
        RECT 1498.780 1593.960 1499.040 1594.220 ;
        RECT 1498.320 1559.620 1498.580 1559.880 ;
        RECT 1498.780 1559.620 1499.040 1559.880 ;
        RECT 1497.860 1511.000 1498.120 1511.260 ;
        RECT 1498.780 1511.000 1499.040 1511.260 ;
        RECT 1498.320 1497.060 1498.580 1497.320 ;
        RECT 1498.780 1449.120 1499.040 1449.380 ;
        RECT 1497.400 1303.940 1497.660 1304.200 ;
        RECT 1498.320 1303.940 1498.580 1304.200 ;
        RECT 1497.400 1159.100 1497.660 1159.360 ;
        RECT 1498.780 1159.100 1499.040 1159.360 ;
        RECT 1497.400 1062.880 1497.660 1063.140 ;
        RECT 1498.780 1062.880 1499.040 1063.140 ;
        RECT 1498.320 1013.920 1498.580 1014.180 ;
        RECT 1498.780 966.320 1499.040 966.580 ;
        RECT 1497.400 869.760 1497.660 870.020 ;
        RECT 1498.780 869.760 1499.040 870.020 ;
        RECT 1497.400 820.800 1497.660 821.060 ;
        RECT 1498.320 820.800 1498.580 821.060 ;
        RECT 1498.320 506.980 1498.580 507.240 ;
        RECT 1498.320 496.440 1498.580 496.700 ;
        RECT 1498.320 434.560 1498.580 434.820 ;
        RECT 1498.320 386.280 1498.580 386.540 ;
        RECT 1498.320 337.660 1498.580 337.920 ;
        RECT 1498.320 304.680 1498.580 304.940 ;
        RECT 406.740 199.280 407.000 199.540 ;
        RECT 1498.780 199.280 1499.040 199.540 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3443.170 1500.820 3517.600 ;
        RECT 1498.320 3442.850 1498.580 3443.170 ;
        RECT 1500.620 3442.850 1500.880 3443.170 ;
        RECT 1498.380 3429.650 1498.520 3442.850 ;
        RECT 1497.920 3429.510 1498.520 3429.650 ;
        RECT 1497.920 3422.430 1498.060 3429.510 ;
        RECT 1497.860 3422.110 1498.120 3422.430 ;
        RECT 1499.700 3332.690 1499.960 3333.010 ;
        RECT 1499.760 3298.410 1499.900 3332.690 ;
        RECT 1498.840 3298.270 1499.900 3298.410 ;
        RECT 1498.840 3236.450 1498.980 3298.270 ;
        RECT 1498.320 3236.130 1498.580 3236.450 ;
        RECT 1498.780 3236.130 1499.040 3236.450 ;
        RECT 1498.380 3202.110 1498.520 3236.130 ;
        RECT 1498.320 3201.790 1498.580 3202.110 ;
        RECT 1498.780 3201.790 1499.040 3202.110 ;
        RECT 1498.840 3153.490 1498.980 3201.790 ;
        RECT 1497.860 3153.170 1498.120 3153.490 ;
        RECT 1498.780 3153.170 1499.040 3153.490 ;
        RECT 1497.920 3152.890 1498.060 3153.170 ;
        RECT 1497.920 3152.750 1498.520 3152.890 ;
        RECT 1498.380 3105.290 1498.520 3152.750 ;
        RECT 1498.380 3105.150 1498.980 3105.290 ;
        RECT 1498.840 3056.930 1498.980 3105.150 ;
        RECT 1497.860 3056.610 1498.120 3056.930 ;
        RECT 1498.780 3056.610 1499.040 3056.930 ;
        RECT 1497.920 3056.330 1498.060 3056.610 ;
        RECT 1497.920 3056.190 1498.520 3056.330 ;
        RECT 1498.380 3042.990 1498.520 3056.190 ;
        RECT 1498.320 3042.670 1498.580 3042.990 ;
        RECT 1499.240 3008.330 1499.500 3008.650 ;
        RECT 1499.300 2994.710 1499.440 3008.330 ;
        RECT 1499.240 2994.390 1499.500 2994.710 ;
        RECT 1499.700 2946.450 1499.960 2946.770 ;
        RECT 1499.760 2912.430 1499.900 2946.450 ;
        RECT 1499.700 2912.110 1499.960 2912.430 ;
        RECT 1499.240 2911.430 1499.500 2911.750 ;
        RECT 1499.300 2863.210 1499.440 2911.430 ;
        RECT 1498.380 2863.070 1499.440 2863.210 ;
        RECT 1498.380 2849.725 1498.520 2863.070 ;
        RECT 1498.310 2849.355 1498.590 2849.725 ;
        RECT 1497.850 2801.755 1498.130 2802.125 ;
        RECT 1497.920 2767.330 1498.060 2801.755 ;
        RECT 1497.920 2767.190 1498.520 2767.330 ;
        RECT 1498.380 2753.310 1498.520 2767.190 ;
        RECT 1497.400 2752.990 1497.660 2753.310 ;
        RECT 1498.320 2752.990 1498.580 2753.310 ;
        RECT 1497.460 2746.365 1497.600 2752.990 ;
        RECT 1496.470 2745.995 1496.750 2746.365 ;
        RECT 1497.390 2745.995 1497.670 2746.365 ;
        RECT 1496.540 2718.630 1496.680 2745.995 ;
        RECT 1496.480 2718.310 1496.740 2718.630 ;
        RECT 1497.400 2718.310 1497.660 2718.630 ;
        RECT 1497.460 2697.970 1497.600 2718.310 ;
        RECT 1497.460 2697.830 1498.060 2697.970 ;
        RECT 1497.920 2656.750 1498.060 2697.830 ;
        RECT 1497.860 2656.430 1498.120 2656.750 ;
        RECT 1498.780 2656.430 1499.040 2656.750 ;
        RECT 1498.840 2622.410 1498.980 2656.430 ;
        RECT 1498.780 2622.090 1499.040 2622.410 ;
        RECT 1499.240 2621.750 1499.500 2622.070 ;
        RECT 1499.300 2608.325 1499.440 2621.750 ;
        RECT 1498.310 2607.955 1498.590 2608.325 ;
        RECT 1499.230 2607.955 1499.510 2608.325 ;
        RECT 1498.380 2560.190 1498.520 2607.955 ;
        RECT 1498.320 2559.870 1498.580 2560.190 ;
        RECT 1499.700 2559.870 1499.960 2560.190 ;
        RECT 1499.760 2511.910 1499.900 2559.870 ;
        RECT 1498.780 2511.765 1499.040 2511.910 ;
        RECT 1497.390 2511.395 1497.670 2511.765 ;
        RECT 1498.770 2511.395 1499.050 2511.765 ;
        RECT 1499.700 2511.590 1499.960 2511.910 ;
        RECT 1497.460 2463.485 1497.600 2511.395 ;
        RECT 1497.390 2463.115 1497.670 2463.485 ;
        RECT 1498.310 2463.115 1498.590 2463.485 ;
        RECT 1498.320 2462.970 1498.580 2463.115 ;
        RECT 1498.320 2428.630 1498.580 2428.950 ;
        RECT 1498.380 2415.090 1498.520 2428.630 ;
        RECT 1498.380 2414.950 1498.980 2415.090 ;
        RECT 1498.840 2380.670 1498.980 2414.950 ;
        RECT 1497.860 2380.410 1498.120 2380.670 ;
        RECT 1497.860 2380.350 1498.520 2380.410 ;
        RECT 1498.780 2380.350 1499.040 2380.670 ;
        RECT 1497.920 2380.270 1498.520 2380.350 ;
        RECT 1498.380 2366.730 1498.520 2380.270 ;
        RECT 1498.320 2366.410 1498.580 2366.730 ;
        RECT 1498.320 2331.730 1498.580 2332.050 ;
        RECT 1498.380 2318.530 1498.520 2331.730 ;
        RECT 1498.380 2318.390 1498.980 2318.530 ;
        RECT 1498.840 2304.510 1498.980 2318.390 ;
        RECT 1496.940 2304.190 1497.200 2304.510 ;
        RECT 1498.780 2304.190 1499.040 2304.510 ;
        RECT 1497.000 2256.650 1497.140 2304.190 ;
        RECT 1497.000 2256.510 1497.600 2256.650 ;
        RECT 1497.460 2249.430 1497.600 2256.510 ;
        RECT 1497.400 2249.110 1497.660 2249.430 ;
        RECT 1497.860 2201.170 1498.120 2201.490 ;
        RECT 1497.920 2184.150 1498.060 2201.170 ;
        RECT 1497.860 2183.830 1498.120 2184.150 ;
        RECT 1497.860 2118.210 1498.120 2118.530 ;
        RECT 1497.920 2111.390 1498.060 2118.210 ;
        RECT 1497.860 2111.070 1498.120 2111.390 ;
        RECT 1498.780 2111.070 1499.040 2111.390 ;
        RECT 1498.840 2063.645 1498.980 2111.070 ;
        RECT 1497.390 2063.275 1497.670 2063.645 ;
        RECT 1498.770 2063.275 1499.050 2063.645 ;
        RECT 1497.460 2063.110 1497.600 2063.275 ;
        RECT 1497.400 2062.790 1497.660 2063.110 ;
        RECT 1497.860 2062.790 1498.120 2063.110 ;
        RECT 1497.920 2008.030 1498.060 2062.790 ;
        RECT 1496.020 2007.710 1496.280 2008.030 ;
        RECT 1497.860 2007.710 1498.120 2008.030 ;
        RECT 1496.080 1960.285 1496.220 2007.710 ;
        RECT 1496.010 1959.915 1496.290 1960.285 ;
        RECT 1496.930 1959.915 1497.210 1960.285 ;
        RECT 1497.000 1959.750 1497.140 1959.915 ;
        RECT 1496.940 1959.430 1497.200 1959.750 ;
        RECT 1497.860 1945.150 1498.120 1945.470 ;
        RECT 1497.920 1897.530 1498.060 1945.150 ;
        RECT 1497.860 1897.210 1498.120 1897.530 ;
        RECT 1498.780 1897.210 1499.040 1897.530 ;
        RECT 1498.840 1859.530 1498.980 1897.210 ;
        RECT 1498.840 1859.390 1499.440 1859.530 ;
        RECT 1499.300 1787.710 1499.440 1859.390 ;
        RECT 1499.240 1787.390 1499.500 1787.710 ;
        RECT 1498.780 1780.650 1499.040 1780.910 ;
        RECT 1498.780 1780.590 1499.440 1780.650 ;
        RECT 1498.840 1780.510 1499.440 1780.590 ;
        RECT 1499.300 1773.430 1499.440 1780.510 ;
        RECT 1499.240 1773.110 1499.500 1773.430 ;
        RECT 1499.700 1683.690 1499.960 1684.010 ;
        RECT 1499.760 1656.890 1499.900 1683.690 ;
        RECT 1499.300 1656.750 1499.900 1656.890 ;
        RECT 1499.300 1635.730 1499.440 1656.750 ;
        RECT 1498.780 1635.410 1499.040 1635.730 ;
        RECT 1499.240 1635.410 1499.500 1635.730 ;
        RECT 1498.840 1594.250 1498.980 1635.410 ;
        RECT 1498.320 1593.930 1498.580 1594.250 ;
        RECT 1498.780 1593.930 1499.040 1594.250 ;
        RECT 1498.380 1559.910 1498.520 1593.930 ;
        RECT 1498.320 1559.590 1498.580 1559.910 ;
        RECT 1498.780 1559.590 1499.040 1559.910 ;
        RECT 1498.840 1511.290 1498.980 1559.590 ;
        RECT 1497.860 1510.970 1498.120 1511.290 ;
        RECT 1498.780 1510.970 1499.040 1511.290 ;
        RECT 1497.920 1510.690 1498.060 1510.970 ;
        RECT 1497.920 1510.550 1498.520 1510.690 ;
        RECT 1498.380 1497.350 1498.520 1510.550 ;
        RECT 1498.320 1497.030 1498.580 1497.350 ;
        RECT 1498.780 1449.090 1499.040 1449.410 ;
        RECT 1498.840 1414.130 1498.980 1449.090 ;
        RECT 1498.380 1413.990 1498.980 1414.130 ;
        RECT 1498.380 1366.645 1498.520 1413.990 ;
        RECT 1498.310 1366.275 1498.590 1366.645 ;
        RECT 1498.310 1352.675 1498.590 1353.045 ;
        RECT 1498.380 1304.230 1498.520 1352.675 ;
        RECT 1497.400 1303.910 1497.660 1304.230 ;
        RECT 1498.320 1303.910 1498.580 1304.230 ;
        RECT 1497.460 1256.485 1497.600 1303.910 ;
        RECT 1497.390 1256.115 1497.670 1256.485 ;
        RECT 1498.770 1256.115 1499.050 1256.485 ;
        RECT 1498.840 1221.010 1498.980 1256.115 ;
        RECT 1498.380 1220.870 1498.980 1221.010 ;
        RECT 1498.380 1207.525 1498.520 1220.870 ;
        RECT 1497.390 1207.155 1497.670 1207.525 ;
        RECT 1498.310 1207.155 1498.590 1207.525 ;
        RECT 1497.460 1159.390 1497.600 1207.155 ;
        RECT 1497.400 1159.070 1497.660 1159.390 ;
        RECT 1498.780 1159.070 1499.040 1159.390 ;
        RECT 1498.840 1124.450 1498.980 1159.070 ;
        RECT 1498.380 1124.310 1498.980 1124.450 ;
        RECT 1498.380 1110.965 1498.520 1124.310 ;
        RECT 1497.390 1110.595 1497.670 1110.965 ;
        RECT 1498.310 1110.595 1498.590 1110.965 ;
        RECT 1497.460 1063.170 1497.600 1110.595 ;
        RECT 1497.400 1062.850 1497.660 1063.170 ;
        RECT 1498.780 1062.850 1499.040 1063.170 ;
        RECT 1498.840 1027.890 1498.980 1062.850 ;
        RECT 1498.380 1027.750 1498.980 1027.890 ;
        RECT 1498.380 1014.210 1498.520 1027.750 ;
        RECT 1498.320 1013.890 1498.580 1014.210 ;
        RECT 1498.780 966.290 1499.040 966.610 ;
        RECT 1498.840 931.330 1498.980 966.290 ;
        RECT 1498.380 931.190 1498.980 931.330 ;
        RECT 1498.380 917.845 1498.520 931.190 ;
        RECT 1497.390 917.475 1497.670 917.845 ;
        RECT 1498.310 917.475 1498.590 917.845 ;
        RECT 1497.460 870.050 1497.600 917.475 ;
        RECT 1497.400 869.730 1497.660 870.050 ;
        RECT 1498.780 869.730 1499.040 870.050 ;
        RECT 1498.840 834.770 1498.980 869.730 ;
        RECT 1498.380 834.630 1498.980 834.770 ;
        RECT 1498.380 821.090 1498.520 834.630 ;
        RECT 1497.400 820.770 1497.660 821.090 ;
        RECT 1498.320 820.770 1498.580 821.090 ;
        RECT 1497.460 773.005 1497.600 820.770 ;
        RECT 1497.390 772.635 1497.670 773.005 ;
        RECT 1498.770 772.635 1499.050 773.005 ;
        RECT 1498.840 738.210 1498.980 772.635 ;
        RECT 1498.380 738.070 1498.980 738.210 ;
        RECT 1498.380 700.130 1498.520 738.070 ;
        RECT 1497.460 699.990 1498.520 700.130 ;
        RECT 1497.460 676.445 1497.600 699.990 ;
        RECT 1497.390 676.075 1497.670 676.445 ;
        RECT 1498.770 676.075 1499.050 676.445 ;
        RECT 1498.840 641.650 1498.980 676.075 ;
        RECT 1498.380 641.510 1498.980 641.650 ;
        RECT 1498.380 603.570 1498.520 641.510 ;
        RECT 1497.460 603.430 1498.520 603.570 ;
        RECT 1497.460 579.885 1497.600 603.430 ;
        RECT 1497.390 579.515 1497.670 579.885 ;
        RECT 1498.770 579.515 1499.050 579.885 ;
        RECT 1498.840 545.090 1498.980 579.515 ;
        RECT 1498.380 544.950 1498.980 545.090 ;
        RECT 1498.380 507.270 1498.520 544.950 ;
        RECT 1498.320 506.950 1498.580 507.270 ;
        RECT 1498.320 496.410 1498.580 496.730 ;
        RECT 1498.380 483.210 1498.520 496.410 ;
        RECT 1498.380 483.070 1498.980 483.210 ;
        RECT 1498.840 448.530 1498.980 483.070 ;
        RECT 1498.380 448.390 1498.980 448.530 ;
        RECT 1498.380 434.850 1498.520 448.390 ;
        RECT 1498.320 434.530 1498.580 434.850 ;
        RECT 1498.320 386.250 1498.580 386.570 ;
        RECT 1498.380 337.950 1498.520 386.250 ;
        RECT 1498.320 337.630 1498.580 337.950 ;
        RECT 1498.320 304.650 1498.580 304.970 ;
        RECT 1498.380 255.410 1498.520 304.650 ;
        RECT 1498.380 255.270 1498.980 255.410 ;
        RECT 406.690 216.000 406.970 220.000 ;
        RECT 406.800 199.570 406.940 216.000 ;
        RECT 1498.840 199.570 1498.980 255.270 ;
        RECT 406.740 199.250 407.000 199.570 ;
        RECT 1498.780 199.250 1499.040 199.570 ;
      LAYER via2 ;
        RECT 1498.310 2849.400 1498.590 2849.680 ;
        RECT 1497.850 2801.800 1498.130 2802.080 ;
        RECT 1496.470 2746.040 1496.750 2746.320 ;
        RECT 1497.390 2746.040 1497.670 2746.320 ;
        RECT 1498.310 2608.000 1498.590 2608.280 ;
        RECT 1499.230 2608.000 1499.510 2608.280 ;
        RECT 1497.390 2511.440 1497.670 2511.720 ;
        RECT 1498.770 2511.440 1499.050 2511.720 ;
        RECT 1497.390 2463.160 1497.670 2463.440 ;
        RECT 1498.310 2463.160 1498.590 2463.440 ;
        RECT 1497.390 2063.320 1497.670 2063.600 ;
        RECT 1498.770 2063.320 1499.050 2063.600 ;
        RECT 1496.010 1959.960 1496.290 1960.240 ;
        RECT 1496.930 1959.960 1497.210 1960.240 ;
        RECT 1498.310 1366.320 1498.590 1366.600 ;
        RECT 1498.310 1352.720 1498.590 1353.000 ;
        RECT 1497.390 1256.160 1497.670 1256.440 ;
        RECT 1498.770 1256.160 1499.050 1256.440 ;
        RECT 1497.390 1207.200 1497.670 1207.480 ;
        RECT 1498.310 1207.200 1498.590 1207.480 ;
        RECT 1497.390 1110.640 1497.670 1110.920 ;
        RECT 1498.310 1110.640 1498.590 1110.920 ;
        RECT 1497.390 917.520 1497.670 917.800 ;
        RECT 1498.310 917.520 1498.590 917.800 ;
        RECT 1497.390 772.680 1497.670 772.960 ;
        RECT 1498.770 772.680 1499.050 772.960 ;
        RECT 1497.390 676.120 1497.670 676.400 ;
        RECT 1498.770 676.120 1499.050 676.400 ;
        RECT 1497.390 579.560 1497.670 579.840 ;
        RECT 1498.770 579.560 1499.050 579.840 ;
      LAYER met3 ;
        RECT 1498.285 2849.700 1498.615 2849.705 ;
        RECT 1498.030 2849.690 1498.615 2849.700 ;
        RECT 1497.830 2849.390 1498.615 2849.690 ;
        RECT 1498.030 2849.380 1498.615 2849.390 ;
        RECT 1498.285 2849.375 1498.615 2849.380 ;
        RECT 1497.825 2802.100 1498.155 2802.105 ;
        RECT 1497.825 2802.090 1498.410 2802.100 ;
        RECT 1497.600 2801.790 1498.410 2802.090 ;
        RECT 1497.825 2801.780 1498.410 2801.790 ;
        RECT 1497.825 2801.775 1498.155 2801.780 ;
        RECT 1496.445 2746.330 1496.775 2746.345 ;
        RECT 1497.365 2746.330 1497.695 2746.345 ;
        RECT 1496.445 2746.030 1497.695 2746.330 ;
        RECT 1496.445 2746.015 1496.775 2746.030 ;
        RECT 1497.365 2746.015 1497.695 2746.030 ;
        RECT 1498.285 2608.290 1498.615 2608.305 ;
        RECT 1499.205 2608.290 1499.535 2608.305 ;
        RECT 1498.285 2607.990 1499.535 2608.290 ;
        RECT 1498.285 2607.975 1498.615 2607.990 ;
        RECT 1499.205 2607.975 1499.535 2607.990 ;
        RECT 1497.365 2511.730 1497.695 2511.745 ;
        RECT 1498.745 2511.730 1499.075 2511.745 ;
        RECT 1497.365 2511.430 1499.075 2511.730 ;
        RECT 1497.365 2511.415 1497.695 2511.430 ;
        RECT 1498.745 2511.415 1499.075 2511.430 ;
        RECT 1497.365 2463.450 1497.695 2463.465 ;
        RECT 1498.285 2463.450 1498.615 2463.465 ;
        RECT 1497.365 2463.150 1498.615 2463.450 ;
        RECT 1497.365 2463.135 1497.695 2463.150 ;
        RECT 1498.285 2463.135 1498.615 2463.150 ;
        RECT 1497.365 2063.610 1497.695 2063.625 ;
        RECT 1498.745 2063.610 1499.075 2063.625 ;
        RECT 1497.365 2063.310 1499.075 2063.610 ;
        RECT 1497.365 2063.295 1497.695 2063.310 ;
        RECT 1498.745 2063.295 1499.075 2063.310 ;
        RECT 1495.985 1960.250 1496.315 1960.265 ;
        RECT 1496.905 1960.250 1497.235 1960.265 ;
        RECT 1495.985 1959.950 1497.235 1960.250 ;
        RECT 1495.985 1959.935 1496.315 1959.950 ;
        RECT 1496.905 1959.935 1497.235 1959.950 ;
        RECT 1498.285 1366.620 1498.615 1366.625 ;
        RECT 1498.030 1366.610 1498.615 1366.620 ;
        RECT 1497.830 1366.310 1498.615 1366.610 ;
        RECT 1498.030 1366.300 1498.615 1366.310 ;
        RECT 1498.285 1366.295 1498.615 1366.300 ;
        RECT 1498.285 1353.020 1498.615 1353.025 ;
        RECT 1498.030 1353.010 1498.615 1353.020 ;
        RECT 1498.030 1352.710 1498.840 1353.010 ;
        RECT 1498.030 1352.700 1498.615 1352.710 ;
        RECT 1498.285 1352.695 1498.615 1352.700 ;
        RECT 1497.365 1256.450 1497.695 1256.465 ;
        RECT 1498.745 1256.450 1499.075 1256.465 ;
        RECT 1497.365 1256.150 1499.075 1256.450 ;
        RECT 1497.365 1256.135 1497.695 1256.150 ;
        RECT 1498.745 1256.135 1499.075 1256.150 ;
        RECT 1497.365 1207.490 1497.695 1207.505 ;
        RECT 1498.285 1207.490 1498.615 1207.505 ;
        RECT 1497.365 1207.190 1498.615 1207.490 ;
        RECT 1497.365 1207.175 1497.695 1207.190 ;
        RECT 1498.285 1207.175 1498.615 1207.190 ;
        RECT 1497.365 1110.930 1497.695 1110.945 ;
        RECT 1498.285 1110.930 1498.615 1110.945 ;
        RECT 1497.365 1110.630 1498.615 1110.930 ;
        RECT 1497.365 1110.615 1497.695 1110.630 ;
        RECT 1498.285 1110.615 1498.615 1110.630 ;
        RECT 1497.365 917.810 1497.695 917.825 ;
        RECT 1498.285 917.810 1498.615 917.825 ;
        RECT 1497.365 917.510 1498.615 917.810 ;
        RECT 1497.365 917.495 1497.695 917.510 ;
        RECT 1498.285 917.495 1498.615 917.510 ;
        RECT 1497.365 772.970 1497.695 772.985 ;
        RECT 1498.745 772.970 1499.075 772.985 ;
        RECT 1497.365 772.670 1499.075 772.970 ;
        RECT 1497.365 772.655 1497.695 772.670 ;
        RECT 1498.745 772.655 1499.075 772.670 ;
        RECT 1497.365 676.410 1497.695 676.425 ;
        RECT 1498.745 676.410 1499.075 676.425 ;
        RECT 1497.365 676.110 1499.075 676.410 ;
        RECT 1497.365 676.095 1497.695 676.110 ;
        RECT 1498.745 676.095 1499.075 676.110 ;
        RECT 1497.365 579.850 1497.695 579.865 ;
        RECT 1498.745 579.850 1499.075 579.865 ;
        RECT 1497.365 579.550 1499.075 579.850 ;
        RECT 1497.365 579.535 1497.695 579.550 ;
        RECT 1498.745 579.535 1499.075 579.550 ;
      LAYER via3 ;
        RECT 1498.060 2849.380 1498.380 2849.700 ;
        RECT 1498.060 2801.780 1498.380 2802.100 ;
        RECT 1498.060 1366.300 1498.380 1366.620 ;
        RECT 1498.060 1352.700 1498.380 1353.020 ;
      LAYER met4 ;
        RECT 1498.055 2849.375 1498.385 2849.705 ;
        RECT 1498.070 2802.105 1498.370 2849.375 ;
        RECT 1498.055 2801.775 1498.385 2802.105 ;
        RECT 1498.055 1366.295 1498.385 1366.625 ;
        RECT 1498.070 1353.025 1498.370 1366.295 ;
        RECT 1498.055 1352.695 1498.385 1353.025 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2038.790 324.260 2039.110 324.320 ;
        RECT 2900.830 324.260 2901.150 324.320 ;
        RECT 2038.790 324.120 2901.150 324.260 ;
        RECT 2038.790 324.060 2039.110 324.120 ;
        RECT 2900.830 324.060 2901.150 324.120 ;
      LAYER via ;
        RECT 2038.820 324.060 2039.080 324.320 ;
        RECT 2900.860 324.060 2901.120 324.320 ;
      LAYER met2 ;
        RECT 512.530 1339.075 512.810 1339.445 ;
        RECT 2038.810 1339.075 2039.090 1339.445 ;
        RECT 512.600 1325.025 512.740 1339.075 ;
        RECT 512.490 1321.025 512.770 1325.025 ;
        RECT 2038.880 324.350 2039.020 1339.075 ;
        RECT 2038.820 324.030 2039.080 324.350 ;
        RECT 2900.860 324.030 2901.120 324.350 ;
        RECT 2900.920 322.845 2901.060 324.030 ;
        RECT 2900.850 322.475 2901.130 322.845 ;
      LAYER via2 ;
        RECT 512.530 1339.120 512.810 1339.400 ;
        RECT 2038.810 1339.120 2039.090 1339.400 ;
        RECT 2900.850 322.520 2901.130 322.800 ;
      LAYER met3 ;
        RECT 512.505 1339.410 512.835 1339.425 ;
        RECT 2038.785 1339.410 2039.115 1339.425 ;
        RECT 512.505 1339.110 2039.115 1339.410 ;
        RECT 512.505 1339.095 512.835 1339.110 ;
        RECT 2038.785 1339.095 2039.115 1339.110 ;
        RECT 2900.825 322.810 2901.155 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2900.825 322.510 2924.800 322.810 ;
        RECT 2900.825 322.495 2901.155 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3503.260 1176.150 3503.320 ;
        RECT 1179.510 3503.260 1179.830 3503.320 ;
        RECT 1175.830 3503.120 1179.830 3503.260 ;
        RECT 1175.830 3503.060 1176.150 3503.120 ;
        RECT 1179.510 3503.060 1179.830 3503.120 ;
        RECT 1179.510 2308.160 1179.830 2308.220 ;
        RECT 1407.670 2308.160 1407.990 2308.220 ;
        RECT 1179.510 2308.020 1407.990 2308.160 ;
        RECT 1179.510 2307.960 1179.830 2308.020 ;
        RECT 1407.670 2307.960 1407.990 2308.020 ;
      LAYER via ;
        RECT 1175.860 3503.060 1176.120 3503.320 ;
        RECT 1179.540 3503.060 1179.800 3503.320 ;
        RECT 1179.540 2307.960 1179.800 2308.220 ;
        RECT 1407.700 2307.960 1407.960 2308.220 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3503.350 1176.060 3517.600 ;
        RECT 1175.860 3503.030 1176.120 3503.350 ;
        RECT 1179.540 3503.030 1179.800 3503.350 ;
        RECT 1179.600 2308.250 1179.740 3503.030 ;
        RECT 1179.540 2307.930 1179.800 2308.250 ;
        RECT 1407.700 2307.930 1407.960 2308.250 ;
        RECT 1407.760 624.765 1407.900 2307.930 ;
        RECT 1407.690 624.395 1407.970 624.765 ;
      LAYER via2 ;
        RECT 1407.690 624.440 1407.970 624.720 ;
      LAYER met3 ;
        RECT 1407.665 624.730 1407.995 624.745 ;
        RECT 1407.665 624.415 1408.210 624.730 ;
        RECT 1407.910 621.920 1408.210 624.415 ;
        RECT 1404.305 621.320 1408.305 621.920 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3502.525 851.760 3517.600 ;
        RECT 851.550 3502.155 851.830 3502.525 ;
        RECT 505.130 216.000 505.410 220.000 ;
        RECT 505.240 205.885 505.380 216.000 ;
        RECT 505.170 205.515 505.450 205.885 ;
      LAYER via2 ;
        RECT 851.550 3502.200 851.830 3502.480 ;
        RECT 505.170 205.560 505.450 205.840 ;
      LAYER met3 ;
        RECT 289.150 3502.490 289.530 3502.500 ;
        RECT 851.525 3502.490 851.855 3502.505 ;
        RECT 289.150 3502.190 851.855 3502.490 ;
        RECT 289.150 3502.180 289.530 3502.190 ;
        RECT 851.525 3502.175 851.855 3502.190 ;
        RECT 289.150 205.850 289.530 205.860 ;
        RECT 505.145 205.850 505.475 205.865 ;
        RECT 289.150 205.550 505.475 205.850 ;
        RECT 289.150 205.540 289.530 205.550 ;
        RECT 505.145 205.535 505.475 205.550 ;
      LAYER via3 ;
        RECT 289.180 3502.180 289.500 3502.500 ;
        RECT 289.180 205.540 289.500 205.860 ;
      LAYER met4 ;
        RECT 289.175 3502.175 289.505 3502.505 ;
        RECT 289.190 205.865 289.490 3502.175 ;
        RECT 289.175 205.535 289.505 205.865 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.230 3503.260 527.550 3503.320 ;
        RECT 848.770 3503.260 849.090 3503.320 ;
        RECT 527.230 3503.120 849.090 3503.260 ;
        RECT 527.230 3503.060 527.550 3503.120 ;
        RECT 848.770 3503.060 849.090 3503.120 ;
      LAYER via ;
        RECT 527.260 3503.060 527.520 3503.320 ;
        RECT 848.800 3503.060 849.060 3503.320 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.350 527.460 3517.600 ;
        RECT 527.260 3503.030 527.520 3503.350 ;
        RECT 848.800 3503.030 849.060 3503.350 ;
        RECT 848.860 1325.730 849.000 3503.030 ;
        RECT 848.860 1325.590 852.220 1325.730 ;
        RECT 852.080 1325.050 852.220 1325.590 ;
        RECT 852.080 1325.025 853.990 1325.050 ;
        RECT 852.080 1324.910 854.090 1325.025 ;
        RECT 853.810 1321.025 854.090 1324.910 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.240 202.790 3502.300 ;
        RECT 206.610 3502.240 206.930 3502.300 ;
        RECT 202.470 3502.100 206.930 3502.240 ;
        RECT 202.470 3502.040 202.790 3502.100 ;
        RECT 206.610 3502.040 206.930 3502.100 ;
        RECT 206.610 211.380 206.930 211.440 ;
        RECT 482.610 211.380 482.930 211.440 ;
        RECT 206.610 211.240 482.930 211.380 ;
        RECT 206.610 211.180 206.930 211.240 ;
        RECT 482.610 211.180 482.930 211.240 ;
        RECT 482.610 206.960 482.930 207.020 ;
        RECT 1083.830 206.960 1084.150 207.020 ;
        RECT 482.610 206.820 1084.150 206.960 ;
        RECT 482.610 206.760 482.930 206.820 ;
        RECT 1083.830 206.760 1084.150 206.820 ;
      LAYER via ;
        RECT 202.500 3502.040 202.760 3502.300 ;
        RECT 206.640 3502.040 206.900 3502.300 ;
        RECT 206.640 211.180 206.900 211.440 ;
        RECT 482.640 211.180 482.900 211.440 ;
        RECT 482.640 206.760 482.900 207.020 ;
        RECT 1083.860 206.760 1084.120 207.020 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.330 202.700 3517.600 ;
        RECT 202.500 3502.010 202.760 3502.330 ;
        RECT 206.640 3502.010 206.900 3502.330 ;
        RECT 206.700 211.470 206.840 3502.010 ;
        RECT 1083.810 216.000 1084.090 220.000 ;
        RECT 206.640 211.150 206.900 211.470 ;
        RECT 482.640 211.150 482.900 211.470 ;
        RECT 482.700 207.050 482.840 211.150 ;
        RECT 1083.920 207.050 1084.060 216.000 ;
        RECT 482.640 206.730 482.900 207.050 ;
        RECT 1083.860 206.730 1084.120 207.050 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 3408.740 16.950 3408.800 ;
        RECT 23.990 3408.740 24.310 3408.800 ;
        RECT 16.630 3408.600 24.310 3408.740 ;
        RECT 16.630 3408.540 16.950 3408.600 ;
        RECT 23.990 3408.540 24.310 3408.600 ;
        RECT 23.990 303.520 24.310 303.580 ;
        RECT 296.770 303.520 297.090 303.580 ;
        RECT 23.990 303.380 297.090 303.520 ;
        RECT 23.990 303.320 24.310 303.380 ;
        RECT 296.770 303.320 297.090 303.380 ;
      LAYER via ;
        RECT 16.660 3408.540 16.920 3408.800 ;
        RECT 24.020 3408.540 24.280 3408.800 ;
        RECT 24.020 303.320 24.280 303.580 ;
        RECT 296.800 303.320 297.060 303.580 ;
      LAYER met2 ;
        RECT 16.650 3411.035 16.930 3411.405 ;
        RECT 16.720 3408.830 16.860 3411.035 ;
        RECT 16.660 3408.510 16.920 3408.830 ;
        RECT 24.020 3408.510 24.280 3408.830 ;
        RECT 24.080 303.610 24.220 3408.510 ;
        RECT 24.020 303.290 24.280 303.610 ;
        RECT 296.800 303.290 297.060 303.610 ;
        RECT 296.860 301.085 297.000 303.290 ;
        RECT 296.790 300.715 297.070 301.085 ;
      LAYER via2 ;
        RECT 16.650 3411.080 16.930 3411.360 ;
        RECT 296.790 300.760 297.070 301.040 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 16.625 3411.370 16.955 3411.385 ;
        RECT -4.800 3411.070 16.955 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 16.625 3411.055 16.955 3411.070 ;
        RECT 296.765 301.050 297.095 301.065 ;
        RECT 296.765 300.960 310.500 301.050 ;
        RECT 296.765 300.750 314.000 300.960 ;
        RECT 296.765 300.735 297.095 300.750 ;
        RECT 310.000 300.360 314.000 300.750 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 3119.060 20.630 3119.120 ;
        RECT 30.890 3119.060 31.210 3119.120 ;
        RECT 20.310 3118.920 31.210 3119.060 ;
        RECT 20.310 3118.860 20.630 3118.920 ;
        RECT 30.890 3118.860 31.210 3118.920 ;
        RECT 30.890 1304.140 31.210 1304.200 ;
        RECT 296.770 1304.140 297.090 1304.200 ;
        RECT 30.890 1304.000 297.090 1304.140 ;
        RECT 30.890 1303.940 31.210 1304.000 ;
        RECT 296.770 1303.940 297.090 1304.000 ;
      LAYER via ;
        RECT 20.340 3118.860 20.600 3119.120 ;
        RECT 30.920 3118.860 31.180 3119.120 ;
        RECT 30.920 1303.940 31.180 1304.200 ;
        RECT 296.800 1303.940 297.060 1304.200 ;
      LAYER met2 ;
        RECT 20.330 3124.075 20.610 3124.445 ;
        RECT 20.400 3119.150 20.540 3124.075 ;
        RECT 20.340 3118.830 20.600 3119.150 ;
        RECT 30.920 3118.830 31.180 3119.150 ;
        RECT 30.980 1304.230 31.120 3118.830 ;
        RECT 30.920 1303.910 31.180 1304.230 ;
        RECT 296.800 1303.910 297.060 1304.230 ;
        RECT 296.860 1302.045 297.000 1303.910 ;
        RECT 296.790 1301.675 297.070 1302.045 ;
      LAYER via2 ;
        RECT 20.330 3124.120 20.610 3124.400 ;
        RECT 296.790 1301.720 297.070 1302.000 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 20.305 3124.410 20.635 3124.425 ;
        RECT -4.800 3124.110 20.635 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 20.305 3124.095 20.635 3124.110 ;
        RECT 296.765 1302.010 297.095 1302.025 ;
        RECT 296.765 1301.920 310.500 1302.010 ;
        RECT 296.765 1301.710 314.000 1301.920 ;
        RECT 296.765 1301.695 297.095 1301.710 ;
        RECT 310.000 1301.320 314.000 1301.710 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 2836.180 20.630 2836.240 ;
        RECT 1276.570 2836.180 1276.890 2836.240 ;
        RECT 20.310 2836.040 1276.890 2836.180 ;
        RECT 20.310 2835.980 20.630 2836.040 ;
        RECT 1276.570 2835.980 1276.890 2836.040 ;
      LAYER via ;
        RECT 20.340 2835.980 20.600 2836.240 ;
        RECT 1276.600 2835.980 1276.860 2836.240 ;
      LAYER met2 ;
        RECT 20.330 2836.435 20.610 2836.805 ;
        RECT 20.400 2836.270 20.540 2836.435 ;
        RECT 20.340 2835.950 20.600 2836.270 ;
        RECT 1276.600 2835.950 1276.860 2836.270 ;
        RECT 1276.660 1325.050 1276.800 2835.950 ;
        RECT 1276.660 1325.025 1279.030 1325.050 ;
        RECT 1276.660 1324.910 1279.130 1325.025 ;
        RECT 1278.850 1321.025 1279.130 1324.910 ;
      LAYER via2 ;
        RECT 20.330 2836.480 20.610 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 20.305 2836.770 20.635 2836.785 ;
        RECT -4.800 2836.470 20.635 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 20.305 2836.455 20.635 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 19.390 2546.500 19.710 2546.560 ;
        RECT 1214.470 2546.500 1214.790 2546.560 ;
        RECT 19.390 2546.360 1214.790 2546.500 ;
        RECT 19.390 2546.300 19.710 2546.360 ;
        RECT 1214.470 2546.300 1214.790 2546.360 ;
      LAYER via ;
        RECT 19.420 2546.300 19.680 2546.560 ;
        RECT 1214.500 2546.300 1214.760 2546.560 ;
      LAYER met2 ;
        RECT 19.410 2549.475 19.690 2549.845 ;
        RECT 19.480 2546.590 19.620 2549.475 ;
        RECT 19.420 2546.270 19.680 2546.590 ;
        RECT 1214.500 2546.270 1214.760 2546.590 ;
        RECT 1214.560 1344.090 1214.700 2546.270 ;
        RECT 1214.560 1343.950 1218.380 1344.090 ;
        RECT 1218.240 1325.050 1218.380 1343.950 ;
        RECT 1218.240 1325.025 1220.150 1325.050 ;
        RECT 1218.240 1324.910 1220.250 1325.025 ;
        RECT 1219.970 1321.025 1220.250 1324.910 ;
      LAYER via2 ;
        RECT 19.410 2549.520 19.690 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 19.385 2549.810 19.715 2549.825 ;
        RECT -4.800 2549.510 19.715 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 19.385 2549.495 19.715 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 217.160 17.410 217.220 ;
        RECT 285.270 217.160 285.590 217.220 ;
        RECT 17.090 217.020 285.590 217.160 ;
        RECT 17.090 216.960 17.410 217.020 ;
        RECT 285.270 216.960 285.590 217.020 ;
        RECT 285.270 205.940 285.590 206.000 ;
        RECT 717.670 205.940 717.990 206.000 ;
        RECT 285.270 205.800 717.990 205.940 ;
        RECT 285.270 205.740 285.590 205.800 ;
        RECT 717.670 205.740 717.990 205.800 ;
      LAYER via ;
        RECT 17.120 216.960 17.380 217.220 ;
        RECT 285.300 216.960 285.560 217.220 ;
        RECT 285.300 205.740 285.560 206.000 ;
        RECT 717.700 205.740 717.960 206.000 ;
      LAYER met2 ;
        RECT 17.110 2261.835 17.390 2262.205 ;
        RECT 17.180 217.250 17.320 2261.835 ;
        RECT 17.120 216.930 17.380 217.250 ;
        RECT 285.300 216.930 285.560 217.250 ;
        RECT 285.360 206.030 285.500 216.930 ;
        RECT 717.650 216.000 717.930 220.000 ;
        RECT 717.760 206.030 717.900 216.000 ;
        RECT 285.300 205.710 285.560 206.030 ;
        RECT 717.700 205.710 717.960 206.030 ;
      LAYER via2 ;
        RECT 17.110 2261.880 17.390 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.085 2262.170 17.415 2262.185 ;
        RECT -4.800 2261.870 17.415 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.085 2261.855 17.415 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 1973.600 20.630 1973.660 ;
        RECT 1408.130 1973.600 1408.450 1973.660 ;
        RECT 20.310 1973.460 1408.450 1973.600 ;
        RECT 20.310 1973.400 20.630 1973.460 ;
        RECT 1408.130 1973.400 1408.450 1973.460 ;
      LAYER via ;
        RECT 20.340 1973.400 20.600 1973.660 ;
        RECT 1408.160 1973.400 1408.420 1973.660 ;
      LAYER met2 ;
        RECT 20.330 1974.875 20.610 1975.245 ;
        RECT 20.400 1973.690 20.540 1974.875 ;
        RECT 20.340 1973.370 20.600 1973.690 ;
        RECT 1408.160 1973.370 1408.420 1973.690 ;
        RECT 1408.220 646.525 1408.360 1973.370 ;
        RECT 1408.150 646.155 1408.430 646.525 ;
      LAYER via2 ;
        RECT 20.330 1974.920 20.610 1975.200 ;
        RECT 1408.150 646.200 1408.430 646.480 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 20.305 1975.210 20.635 1975.225 ;
        RECT -4.800 1974.910 20.635 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 20.305 1974.895 20.635 1974.910 ;
        RECT 1408.125 646.490 1408.455 646.505 ;
        RECT 1407.910 646.175 1408.455 646.490 ;
        RECT 1407.910 643.680 1408.210 646.175 ;
        RECT 1404.305 643.080 1408.305 643.680 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 665.195 301.210 665.565 ;
        RECT 301.000 407.845 301.140 665.195 ;
        RECT 300.930 407.475 301.210 407.845 ;
      LAYER via2 ;
        RECT 300.930 665.240 301.210 665.520 ;
        RECT 300.930 407.520 301.210 407.800 ;
      LAYER met3 ;
        RECT 300.905 665.530 301.235 665.545 ;
        RECT 300.905 665.440 310.500 665.530 ;
        RECT 300.905 665.230 314.000 665.440 ;
        RECT 300.905 665.215 301.235 665.230 ;
        RECT 310.000 664.840 314.000 665.230 ;
        RECT 2901.950 557.410 2902.330 557.420 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2901.950 557.110 2924.800 557.410 ;
        RECT 2901.950 557.100 2902.330 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 300.905 407.810 301.235 407.825 ;
        RECT 305.710 407.810 306.090 407.820 ;
        RECT 300.905 407.510 306.090 407.810 ;
        RECT 300.905 407.495 301.235 407.510 ;
        RECT 305.710 407.500 306.090 407.510 ;
        RECT 1441.910 365.650 1442.290 365.660 ;
        RECT 1489.750 365.650 1490.130 365.660 ;
        RECT 1441.910 365.350 1490.130 365.650 ;
        RECT 1441.910 365.340 1442.290 365.350 ;
        RECT 1489.750 365.340 1490.130 365.350 ;
        RECT 2763.030 365.650 2763.410 365.660 ;
        RECT 2767.630 365.650 2768.010 365.660 ;
        RECT 2763.030 365.350 2768.010 365.650 ;
        RECT 2763.030 365.340 2763.410 365.350 ;
        RECT 2767.630 365.340 2768.010 365.350 ;
        RECT 1406.950 362.250 1407.330 362.260 ;
        RECT 1417.070 362.250 1417.450 362.260 ;
        RECT 1406.950 361.950 1417.450 362.250 ;
        RECT 1406.950 361.940 1407.330 361.950 ;
        RECT 1417.070 361.940 1417.450 361.950 ;
        RECT 1892.710 362.250 1893.090 362.260 ;
        RECT 1931.350 362.250 1931.730 362.260 ;
        RECT 1892.710 361.950 1931.730 362.250 ;
        RECT 1892.710 361.940 1893.090 361.950 ;
        RECT 1931.350 361.940 1931.730 361.950 ;
        RECT 2078.550 362.250 2078.930 362.260 ;
        RECT 2124.550 362.250 2124.930 362.260 ;
        RECT 2078.550 361.950 2124.930 362.250 ;
        RECT 2078.550 361.940 2078.930 361.950 ;
        RECT 2124.550 361.940 2124.930 361.950 ;
        RECT 2186.190 362.250 2186.570 362.260 ;
        RECT 2221.150 362.250 2221.530 362.260 ;
        RECT 2186.190 361.950 2221.530 362.250 ;
        RECT 2186.190 361.940 2186.570 361.950 ;
        RECT 2221.150 361.940 2221.530 361.950 ;
        RECT 2376.630 362.250 2377.010 362.260 ;
        RECT 2381.230 362.250 2381.610 362.260 ;
        RECT 2376.630 361.950 2381.610 362.250 ;
        RECT 2376.630 361.940 2377.010 361.950 ;
        RECT 2381.230 361.940 2381.610 361.950 ;
        RECT 1545.870 358.850 1546.250 358.860 ;
        RECT 1592.790 358.850 1593.170 358.860 ;
        RECT 1545.870 358.550 1593.170 358.850 ;
        RECT 1545.870 358.540 1546.250 358.550 ;
        RECT 1592.790 358.540 1593.170 358.550 ;
        RECT 1642.470 358.850 1642.850 358.860 ;
        RECT 1689.390 358.850 1689.770 358.860 ;
        RECT 1642.470 358.550 1689.770 358.850 ;
        RECT 1642.470 358.540 1642.850 358.550 ;
        RECT 1689.390 358.540 1689.770 358.550 ;
        RECT 1739.070 358.850 1739.450 358.860 ;
        RECT 1785.990 358.850 1786.370 358.860 ;
        RECT 1739.070 358.550 1786.370 358.850 ;
        RECT 1739.070 358.540 1739.450 358.550 ;
        RECT 1785.990 358.540 1786.370 358.550 ;
        RECT 1835.670 358.850 1836.050 358.860 ;
        RECT 1882.590 358.850 1882.970 358.860 ;
        RECT 1835.670 358.550 1882.970 358.850 ;
        RECT 1835.670 358.540 1836.050 358.550 ;
        RECT 1882.590 358.540 1882.970 358.550 ;
        RECT 2269.910 358.850 2270.290 358.860 ;
        RECT 2317.750 358.850 2318.130 358.860 ;
        RECT 2269.910 358.550 2318.130 358.850 ;
        RECT 2269.910 358.540 2270.290 358.550 ;
        RECT 2317.750 358.540 2318.130 358.550 ;
        RECT 2511.870 358.850 2512.250 358.860 ;
        RECT 2558.790 358.850 2559.170 358.860 ;
        RECT 2511.870 358.550 2559.170 358.850 ;
        RECT 2511.870 358.540 2512.250 358.550 ;
        RECT 2558.790 358.540 2559.170 358.550 ;
      LAYER via3 ;
        RECT 2901.980 557.100 2902.300 557.420 ;
        RECT 305.740 407.500 306.060 407.820 ;
        RECT 1441.940 365.340 1442.260 365.660 ;
        RECT 1489.780 365.340 1490.100 365.660 ;
        RECT 2763.060 365.340 2763.380 365.660 ;
        RECT 2767.660 365.340 2767.980 365.660 ;
        RECT 1406.980 361.940 1407.300 362.260 ;
        RECT 1417.100 361.940 1417.420 362.260 ;
        RECT 1892.740 361.940 1893.060 362.260 ;
        RECT 1931.380 361.940 1931.700 362.260 ;
        RECT 2078.580 361.940 2078.900 362.260 ;
        RECT 2124.580 361.940 2124.900 362.260 ;
        RECT 2186.220 361.940 2186.540 362.260 ;
        RECT 2221.180 361.940 2221.500 362.260 ;
        RECT 2376.660 361.940 2376.980 362.260 ;
        RECT 2381.260 361.940 2381.580 362.260 ;
        RECT 1545.900 358.540 1546.220 358.860 ;
        RECT 1592.820 358.540 1593.140 358.860 ;
        RECT 1642.500 358.540 1642.820 358.860 ;
        RECT 1689.420 358.540 1689.740 358.860 ;
        RECT 1739.100 358.540 1739.420 358.860 ;
        RECT 1786.020 358.540 1786.340 358.860 ;
        RECT 1835.700 358.540 1836.020 358.860 ;
        RECT 1882.620 358.540 1882.940 358.860 ;
        RECT 2269.940 358.540 2270.260 358.860 ;
        RECT 2317.780 358.540 2318.100 358.860 ;
        RECT 2511.900 358.540 2512.220 358.860 ;
        RECT 2558.820 358.540 2559.140 358.860 ;
      LAYER met4 ;
        RECT 2901.975 557.095 2902.305 557.425 ;
        RECT 305.735 407.495 306.065 407.825 ;
        RECT 305.750 362.690 306.050 407.495 ;
        RECT 2901.990 366.090 2902.290 557.095 ;
        RECT 1416.670 364.910 1417.850 366.090 ;
        RECT 1441.510 364.910 1442.690 366.090 ;
        RECT 1489.350 364.910 1490.530 366.090 ;
        RECT 1930.950 364.910 1932.130 366.090 ;
        RECT 2762.630 364.910 2763.810 366.090 ;
        RECT 2767.230 364.910 2768.410 366.090 ;
        RECT 2901.550 364.910 2902.730 366.090 ;
        RECT 305.310 361.510 306.490 362.690 ;
        RECT 1406.550 361.510 1407.730 362.690 ;
        RECT 1417.110 362.265 1417.410 364.910 ;
        RECT 1417.095 361.935 1417.425 362.265 ;
        RECT 1592.390 361.510 1593.570 362.690 ;
        RECT 1688.990 361.510 1690.170 362.690 ;
        RECT 1785.590 361.510 1786.770 362.690 ;
        RECT 1882.190 361.510 1883.370 362.690 ;
        RECT 1892.310 361.510 1893.490 362.690 ;
        RECT 1931.390 362.265 1931.690 364.910 ;
        RECT 1931.375 361.935 1931.705 362.265 ;
        RECT 2078.150 361.510 2079.330 362.690 ;
        RECT 2124.575 361.935 2124.905 362.265 ;
        RECT 1545.470 358.110 1546.650 359.290 ;
        RECT 1592.830 358.865 1593.130 361.510 ;
        RECT 1592.815 358.535 1593.145 358.865 ;
        RECT 1642.070 358.110 1643.250 359.290 ;
        RECT 1689.430 358.865 1689.730 361.510 ;
        RECT 1689.415 358.535 1689.745 358.865 ;
        RECT 1738.670 358.110 1739.850 359.290 ;
        RECT 1786.030 358.865 1786.330 361.510 ;
        RECT 1786.015 358.535 1786.345 358.865 ;
        RECT 1835.270 358.110 1836.450 359.290 ;
        RECT 1882.630 358.865 1882.930 361.510 ;
        RECT 2124.590 359.290 2124.890 361.935 ;
        RECT 2185.790 361.510 2186.970 362.690 ;
        RECT 2220.750 361.510 2221.930 362.690 ;
        RECT 2376.230 361.510 2377.410 362.690 ;
        RECT 2380.830 361.510 2382.010 362.690 ;
        RECT 1882.615 358.535 1882.945 358.865 ;
        RECT 2028.470 358.110 2029.650 359.290 ;
        RECT 2124.150 358.110 2125.330 359.290 ;
        RECT 2269.510 358.110 2270.690 359.290 ;
        RECT 2317.350 358.110 2318.530 359.290 ;
        RECT 2511.470 358.110 2512.650 359.290 ;
        RECT 2558.390 358.110 2559.570 359.290 ;
        RECT 2028.910 349.090 2029.210 358.110 ;
        RECT 2028.470 347.910 2029.650 349.090 ;
      LAYER met5 ;
        RECT 349.260 364.700 436.420 366.300 ;
        RECT 349.260 362.900 350.860 364.700 ;
        RECT 305.100 361.300 350.860 362.900 ;
        RECT 398.940 357.900 401.460 364.700 ;
        RECT 434.820 359.500 436.420 364.700 ;
        RECT 497.380 364.700 533.020 366.300 ;
        RECT 497.380 359.500 498.980 364.700 ;
        RECT 434.820 357.900 437.340 359.500 ;
        RECT 435.740 345.900 437.340 357.900 ;
        RECT 480.820 357.900 498.980 359.500 ;
        RECT 531.420 359.500 533.020 364.700 ;
        RECT 593.980 364.700 629.620 366.300 ;
        RECT 593.980 359.500 595.580 364.700 ;
        RECT 531.420 357.900 533.940 359.500 ;
        RECT 480.820 345.900 482.420 357.900 ;
        RECT 435.740 344.300 482.420 345.900 ;
        RECT 532.340 345.900 533.940 357.900 ;
        RECT 577.420 357.900 595.580 359.500 ;
        RECT 628.020 359.500 629.620 364.700 ;
        RECT 690.580 364.700 726.220 366.300 ;
        RECT 690.580 359.500 692.180 364.700 ;
        RECT 628.020 357.900 630.540 359.500 ;
        RECT 577.420 345.900 579.020 357.900 ;
        RECT 532.340 344.300 579.020 345.900 ;
        RECT 628.940 345.900 630.540 357.900 ;
        RECT 674.020 357.900 692.180 359.500 ;
        RECT 724.620 359.500 726.220 364.700 ;
        RECT 787.180 364.700 822.820 366.300 ;
        RECT 787.180 359.500 788.780 364.700 ;
        RECT 724.620 357.900 727.140 359.500 ;
        RECT 674.020 345.900 675.620 357.900 ;
        RECT 628.940 344.300 675.620 345.900 ;
        RECT 725.540 345.900 727.140 357.900 ;
        RECT 770.620 357.900 788.780 359.500 ;
        RECT 821.220 359.500 822.820 364.700 ;
        RECT 883.780 364.700 919.420 366.300 ;
        RECT 883.780 359.500 885.380 364.700 ;
        RECT 821.220 357.900 823.740 359.500 ;
        RECT 770.620 345.900 772.220 357.900 ;
        RECT 725.540 344.300 772.220 345.900 ;
        RECT 822.140 345.900 823.740 357.900 ;
        RECT 867.220 357.900 885.380 359.500 ;
        RECT 917.820 359.500 919.420 364.700 ;
        RECT 980.380 364.700 1016.020 366.300 ;
        RECT 980.380 359.500 981.980 364.700 ;
        RECT 917.820 357.900 920.340 359.500 ;
        RECT 867.220 345.900 868.820 357.900 ;
        RECT 822.140 344.300 868.820 345.900 ;
        RECT 918.740 345.900 920.340 357.900 ;
        RECT 963.820 357.900 981.980 359.500 ;
        RECT 1014.420 359.500 1016.020 364.700 ;
        RECT 1076.980 364.700 1112.620 366.300 ;
        RECT 1076.980 359.500 1078.580 364.700 ;
        RECT 1014.420 357.900 1016.940 359.500 ;
        RECT 963.820 345.900 965.420 357.900 ;
        RECT 918.740 344.300 965.420 345.900 ;
        RECT 1015.340 345.900 1016.940 357.900 ;
        RECT 1060.420 357.900 1078.580 359.500 ;
        RECT 1111.020 359.500 1112.620 364.700 ;
        RECT 1173.580 364.700 1209.220 366.300 ;
        RECT 1173.580 359.500 1175.180 364.700 ;
        RECT 1111.020 357.900 1113.540 359.500 ;
        RECT 1060.420 345.900 1062.020 357.900 ;
        RECT 1015.340 344.300 1062.020 345.900 ;
        RECT 1111.940 345.900 1113.540 357.900 ;
        RECT 1157.020 357.900 1175.180 359.500 ;
        RECT 1207.620 359.500 1209.220 364.700 ;
        RECT 1270.180 364.700 1328.820 366.300 ;
        RECT 1416.460 364.700 1442.900 366.300 ;
        RECT 1489.140 364.700 1498.100 366.300 ;
        RECT 1930.740 364.700 1946.140 366.300 ;
        RECT 1270.180 359.500 1271.780 364.700 ;
        RECT 1207.620 357.900 1210.140 359.500 ;
        RECT 1157.020 345.900 1158.620 357.900 ;
        RECT 1111.940 344.300 1158.620 345.900 ;
        RECT 1208.540 345.900 1210.140 357.900 ;
        RECT 1253.620 357.900 1271.780 359.500 ;
        RECT 1327.220 359.500 1328.820 364.700 ;
        RECT 1496.500 362.900 1498.100 364.700 ;
        RECT 1365.860 361.300 1407.940 362.900 ;
        RECT 1496.500 361.300 1545.940 362.900 ;
        RECT 1592.180 361.300 1607.580 362.900 ;
        RECT 1688.780 361.300 1704.180 362.900 ;
        RECT 1785.380 361.300 1800.780 362.900 ;
        RECT 1881.980 361.300 1893.700 362.900 ;
        RECT 1365.860 359.500 1367.460 361.300 ;
        RECT 1327.220 357.900 1367.460 359.500 ;
        RECT 1544.340 359.500 1545.940 361.300 ;
        RECT 1605.980 359.500 1607.580 361.300 ;
        RECT 1702.580 359.500 1704.180 361.300 ;
        RECT 1799.180 359.500 1800.780 361.300 ;
        RECT 1944.540 359.500 1946.140 364.700 ;
        RECT 2571.980 364.700 2643.500 366.300 ;
        RECT 1948.220 361.300 1992.140 362.900 ;
        RECT 1948.220 359.500 1949.820 361.300 ;
        RECT 1544.340 357.900 1546.860 359.500 ;
        RECT 1605.980 357.900 1643.460 359.500 ;
        RECT 1702.580 357.900 1740.060 359.500 ;
        RECT 1799.180 357.900 1836.660 359.500 ;
        RECT 1944.540 357.900 1949.820 359.500 ;
        RECT 1990.540 359.500 1992.140 361.300 ;
        RECT 2074.260 361.300 2079.540 362.900 ;
        RECT 2124.860 361.300 2187.180 362.900 ;
        RECT 2220.540 361.300 2223.980 362.900 ;
        RECT 1990.540 357.900 2029.860 359.500 ;
        RECT 1253.620 345.900 1255.220 357.900 ;
        RECT 2074.260 349.300 2075.860 361.300 ;
        RECT 2124.860 359.500 2126.460 361.300 ;
        RECT 2123.160 357.900 2126.460 359.500 ;
        RECT 2222.380 359.500 2223.980 361.300 ;
        RECT 2364.980 361.300 2377.620 362.900 ;
        RECT 2380.620 361.300 2426.380 362.900 ;
        RECT 2364.980 359.500 2366.580 361.300 ;
        RECT 2222.380 357.900 2270.900 359.500 ;
        RECT 2317.140 357.900 2366.580 359.500 ;
        RECT 2424.780 359.500 2426.380 361.300 ;
        RECT 2431.220 361.300 2475.140 362.900 ;
        RECT 2431.220 359.500 2432.820 361.300 ;
        RECT 2424.780 357.900 2432.820 359.500 ;
        RECT 2473.540 359.500 2475.140 361.300 ;
        RECT 2571.980 359.500 2573.580 364.700 ;
        RECT 2473.540 357.900 2512.860 359.500 ;
        RECT 2558.180 357.900 2573.580 359.500 ;
        RECT 2641.900 359.500 2643.500 364.700 ;
        RECT 2672.260 364.700 2764.020 366.300 ;
        RECT 2767.020 364.700 2815.540 366.300 ;
        RECT 2672.260 359.500 2673.860 364.700 ;
        RECT 2641.900 357.900 2673.860 359.500 ;
        RECT 2813.940 359.500 2815.540 364.700 ;
        RECT 2834.180 364.700 2902.940 366.300 ;
        RECT 2834.180 359.500 2835.780 364.700 ;
        RECT 2813.940 357.900 2835.780 359.500 ;
        RECT 2028.260 347.700 2075.860 349.300 ;
        RECT 1208.540 344.300 1255.220 345.900 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 1683.920 20.630 1683.980 ;
        RECT 1409.510 1683.920 1409.830 1683.980 ;
        RECT 20.310 1683.780 1409.830 1683.920 ;
        RECT 20.310 1683.720 20.630 1683.780 ;
        RECT 1409.510 1683.720 1409.830 1683.780 ;
      LAYER via ;
        RECT 20.340 1683.720 20.600 1683.980 ;
        RECT 1409.540 1683.720 1409.800 1683.980 ;
      LAYER met2 ;
        RECT 20.330 1687.235 20.610 1687.605 ;
        RECT 20.400 1684.010 20.540 1687.235 ;
        RECT 20.340 1683.690 20.600 1684.010 ;
        RECT 1409.540 1683.690 1409.800 1684.010 ;
        RECT 1409.600 418.045 1409.740 1683.690 ;
        RECT 1409.530 417.675 1409.810 418.045 ;
      LAYER via2 ;
        RECT 20.330 1687.280 20.610 1687.560 ;
        RECT 1409.530 417.720 1409.810 418.000 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 20.305 1687.570 20.635 1687.585 ;
        RECT -4.800 1687.270 20.635 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 20.305 1687.255 20.635 1687.270 ;
        RECT 1409.505 418.010 1409.835 418.025 ;
        RECT 1408.060 417.920 1409.835 418.010 ;
        RECT 1404.305 417.710 1409.835 417.920 ;
        RECT 1404.305 417.320 1408.305 417.710 ;
        RECT 1409.505 417.695 1409.835 417.710 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1470.060 16.030 1470.120 ;
        RECT 37.790 1470.060 38.110 1470.120 ;
        RECT 15.710 1469.920 38.110 1470.060 ;
        RECT 15.710 1469.860 16.030 1469.920 ;
        RECT 37.790 1469.860 38.110 1469.920 ;
        RECT 37.790 206.620 38.110 206.680 ;
        RECT 638.550 206.620 638.870 206.680 ;
        RECT 37.790 206.480 638.870 206.620 ;
        RECT 37.790 206.420 38.110 206.480 ;
        RECT 638.550 206.420 638.870 206.480 ;
      LAYER via ;
        RECT 15.740 1469.860 16.000 1470.120 ;
        RECT 37.820 1469.860 38.080 1470.120 ;
        RECT 37.820 206.420 38.080 206.680 ;
        RECT 638.580 206.420 638.840 206.680 ;
      LAYER met2 ;
        RECT 15.730 1471.675 16.010 1472.045 ;
        RECT 15.800 1470.150 15.940 1471.675 ;
        RECT 15.740 1469.830 16.000 1470.150 ;
        RECT 37.820 1469.830 38.080 1470.150 ;
        RECT 37.880 206.710 38.020 1469.830 ;
        RECT 638.530 216.000 638.810 220.000 ;
        RECT 638.640 206.710 638.780 216.000 ;
        RECT 37.820 206.390 38.080 206.710 ;
        RECT 638.580 206.390 638.840 206.710 ;
      LAYER via2 ;
        RECT 15.730 1471.720 16.010 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 15.705 1472.010 16.035 1472.025 ;
        RECT -4.800 1471.710 16.035 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 15.705 1471.695 16.035 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 1256.200 20.630 1256.260 ;
        RECT 44.690 1256.200 45.010 1256.260 ;
        RECT 20.310 1256.060 45.010 1256.200 ;
        RECT 20.310 1256.000 20.630 1256.060 ;
        RECT 44.690 1256.000 45.010 1256.060 ;
        RECT 44.690 206.960 45.010 207.020 ;
        RECT 440.750 206.960 441.070 207.020 ;
        RECT 44.690 206.820 441.070 206.960 ;
        RECT 44.690 206.760 45.010 206.820 ;
        RECT 440.750 206.760 441.070 206.820 ;
      LAYER via ;
        RECT 20.340 1256.000 20.600 1256.260 ;
        RECT 44.720 1256.000 44.980 1256.260 ;
        RECT 44.720 206.760 44.980 207.020 ;
        RECT 440.780 206.760 441.040 207.020 ;
      LAYER met2 ;
        RECT 20.330 1256.115 20.610 1256.485 ;
        RECT 20.340 1255.970 20.600 1256.115 ;
        RECT 44.720 1255.970 44.980 1256.290 ;
        RECT 44.780 207.050 44.920 1255.970 ;
        RECT 440.730 216.000 441.010 220.000 ;
        RECT 440.840 207.050 440.980 216.000 ;
        RECT 44.720 206.730 44.980 207.050 ;
        RECT 440.780 206.730 441.040 207.050 ;
      LAYER via2 ;
        RECT 20.330 1256.160 20.610 1256.440 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 20.305 1256.450 20.635 1256.465 ;
        RECT -4.800 1256.150 20.635 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 20.305 1256.135 20.635 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.810 1207.155 1418.090 1207.525 ;
        RECT 1417.880 1159.925 1418.020 1207.155 ;
        RECT 1417.810 1159.555 1418.090 1159.925 ;
        RECT 1419.190 962.355 1419.470 962.725 ;
        RECT 1419.260 902.205 1419.400 962.355 ;
        RECT 1419.190 901.835 1419.470 902.205 ;
      LAYER via2 ;
        RECT 1417.810 1207.200 1418.090 1207.480 ;
        RECT 1417.810 1159.600 1418.090 1159.880 ;
        RECT 1419.190 962.400 1419.470 962.680 ;
        RECT 1419.190 901.880 1419.470 902.160 ;
      LAYER met3 ;
        RECT 1410.630 1242.170 1411.010 1242.180 ;
        RECT 1417.990 1242.170 1418.370 1242.180 ;
        RECT 1410.630 1241.870 1418.370 1242.170 ;
        RECT 1410.630 1241.860 1411.010 1241.870 ;
        RECT 1417.990 1241.860 1418.370 1241.870 ;
        RECT 1416.150 1221.090 1416.530 1221.100 ;
        RECT 1417.990 1221.090 1418.370 1221.100 ;
        RECT 1416.150 1220.790 1418.370 1221.090 ;
        RECT 1416.150 1220.780 1416.530 1220.790 ;
        RECT 1417.990 1220.780 1418.370 1220.790 ;
        RECT 1416.150 1207.490 1416.530 1207.500 ;
        RECT 1417.785 1207.490 1418.115 1207.505 ;
        RECT 1416.150 1207.190 1418.115 1207.490 ;
        RECT 1416.150 1207.180 1416.530 1207.190 ;
        RECT 1417.785 1207.175 1418.115 1207.190 ;
        RECT 1417.785 1159.900 1418.115 1159.905 ;
        RECT 1417.785 1159.890 1418.370 1159.900 ;
        RECT 1417.560 1159.590 1418.370 1159.890 ;
        RECT 1417.785 1159.580 1418.370 1159.590 ;
        RECT 1417.785 1159.575 1418.115 1159.580 ;
        RECT 1416.150 1100.730 1416.530 1100.740 ;
        RECT 1417.990 1100.730 1418.370 1100.740 ;
        RECT 1416.150 1100.430 1418.370 1100.730 ;
        RECT 1416.150 1100.420 1416.530 1100.430 ;
        RECT 1417.990 1100.420 1418.370 1100.430 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 3.070 1041.270 305.130 1041.570 ;
        RECT 3.070 1040.890 3.370 1041.270 ;
        RECT -4.800 1040.590 3.370 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 304.830 1040.210 305.130 1041.270 ;
        RECT 308.470 1040.210 308.850 1040.220 ;
        RECT 304.830 1039.910 308.850 1040.210 ;
        RECT 308.470 1039.900 308.850 1039.910 ;
        RECT 1416.150 1031.370 1416.530 1031.380 ;
        RECT 1419.830 1031.370 1420.210 1031.380 ;
        RECT 1416.150 1031.070 1420.210 1031.370 ;
        RECT 1416.150 1031.060 1416.530 1031.070 ;
        RECT 1419.830 1031.060 1420.210 1031.070 ;
        RECT 1419.165 962.690 1419.495 962.705 ;
        RECT 1419.830 962.690 1420.210 962.700 ;
        RECT 1419.165 962.390 1420.210 962.690 ;
        RECT 1419.165 962.375 1419.495 962.390 ;
        RECT 1419.830 962.380 1420.210 962.390 ;
        RECT 1416.150 902.170 1416.530 902.180 ;
        RECT 1419.165 902.170 1419.495 902.185 ;
        RECT 1416.150 901.870 1419.495 902.170 ;
        RECT 1416.150 901.860 1416.530 901.870 ;
        RECT 1419.165 901.855 1419.495 901.870 ;
        RECT 1416.150 872.930 1416.530 872.940 ;
        RECT 1418.910 872.930 1419.290 872.940 ;
        RECT 1416.150 872.630 1419.290 872.930 ;
        RECT 1416.150 872.620 1416.530 872.630 ;
        RECT 1418.910 872.620 1419.290 872.630 ;
        RECT 1418.910 812.410 1419.290 812.420 ;
        RECT 1408.060 812.320 1419.290 812.410 ;
        RECT 1404.305 812.110 1419.290 812.320 ;
        RECT 1404.305 811.720 1408.305 812.110 ;
        RECT 1418.910 812.100 1419.290 812.110 ;
      LAYER via3 ;
        RECT 1410.660 1241.860 1410.980 1242.180 ;
        RECT 1418.020 1241.860 1418.340 1242.180 ;
        RECT 1416.180 1220.780 1416.500 1221.100 ;
        RECT 1418.020 1220.780 1418.340 1221.100 ;
        RECT 1416.180 1207.180 1416.500 1207.500 ;
        RECT 1418.020 1159.580 1418.340 1159.900 ;
        RECT 1416.180 1100.420 1416.500 1100.740 ;
        RECT 1418.020 1100.420 1418.340 1100.740 ;
        RECT 308.500 1039.900 308.820 1040.220 ;
        RECT 1416.180 1031.060 1416.500 1031.380 ;
        RECT 1419.860 1031.060 1420.180 1031.380 ;
        RECT 1419.860 962.380 1420.180 962.700 ;
        RECT 1416.180 901.860 1416.500 902.180 ;
        RECT 1416.180 872.620 1416.500 872.940 ;
        RECT 1418.940 872.620 1419.260 872.940 ;
        RECT 1418.940 812.100 1419.260 812.420 ;
      LAYER met4 ;
        RECT 308.070 1242.110 309.250 1243.290 ;
        RECT 1410.230 1242.110 1411.410 1243.290 ;
        RECT 308.510 1040.225 308.810 1242.110 ;
        RECT 1410.655 1241.855 1410.985 1242.110 ;
        RECT 1418.015 1241.855 1418.345 1242.185 ;
        RECT 1418.030 1221.105 1418.330 1241.855 ;
        RECT 1416.175 1220.775 1416.505 1221.105 ;
        RECT 1418.015 1220.775 1418.345 1221.105 ;
        RECT 1416.190 1207.505 1416.490 1220.775 ;
        RECT 1416.175 1207.175 1416.505 1207.505 ;
        RECT 1418.015 1159.575 1418.345 1159.905 ;
        RECT 1418.030 1100.745 1418.330 1159.575 ;
        RECT 1416.175 1100.415 1416.505 1100.745 ;
        RECT 1418.015 1100.415 1418.345 1100.745 ;
        RECT 308.495 1039.895 308.825 1040.225 ;
        RECT 1416.190 1031.385 1416.490 1100.415 ;
        RECT 1416.175 1031.055 1416.505 1031.385 ;
        RECT 1419.855 1031.055 1420.185 1031.385 ;
        RECT 1419.870 962.705 1420.170 1031.055 ;
        RECT 1419.855 962.375 1420.185 962.705 ;
        RECT 1416.175 901.855 1416.505 902.185 ;
        RECT 1416.190 872.945 1416.490 901.855 ;
        RECT 1416.175 872.615 1416.505 872.945 ;
        RECT 1418.935 872.615 1419.265 872.945 ;
        RECT 1418.950 812.425 1419.250 872.615 ;
        RECT 1418.935 812.095 1419.265 812.425 ;
      LAYER via4 ;
        RECT 1410.230 1242.110 1411.410 1243.290 ;
      LAYER met5 ;
        RECT 405.380 1252.100 412.500 1253.700 ;
        RECT 388.820 1248.700 395.940 1250.300 ;
        RECT 388.820 1243.500 390.420 1248.700 ;
        RECT 394.340 1246.900 395.940 1248.700 ;
        RECT 405.380 1246.900 406.980 1252.100 ;
        RECT 394.340 1245.300 406.980 1246.900 ;
        RECT 410.900 1246.900 412.500 1252.100 ;
        RECT 501.060 1248.700 506.340 1250.300 ;
        RECT 410.900 1245.300 420.780 1246.900 ;
        RECT 307.860 1241.900 390.420 1243.500 ;
        RECT 419.180 1243.500 420.780 1245.300 ;
        RECT 501.060 1243.500 502.660 1248.700 ;
        RECT 504.740 1246.900 506.340 1248.700 ;
        RECT 512.100 1248.700 518.300 1250.300 ;
        RECT 512.100 1246.900 513.700 1248.700 ;
        RECT 504.740 1245.300 513.700 1246.900 ;
        RECT 419.180 1241.900 502.660 1243.500 ;
        RECT 516.700 1243.500 518.300 1248.700 ;
        RECT 534.180 1248.700 554.180 1250.300 ;
        RECT 534.180 1243.500 535.780 1248.700 ;
        RECT 516.700 1241.900 535.780 1243.500 ;
        RECT 552.580 1243.500 554.180 1248.700 ;
        RECT 605.940 1245.300 624.100 1246.900 ;
        RECT 605.940 1243.500 607.540 1245.300 ;
        RECT 552.580 1241.900 607.540 1243.500 ;
        RECT 622.500 1243.500 624.100 1245.300 ;
        RECT 702.540 1245.300 721.620 1246.900 ;
        RECT 702.540 1243.500 704.140 1245.300 ;
        RECT 622.500 1241.900 704.140 1243.500 ;
        RECT 720.020 1243.500 721.620 1245.300 ;
        RECT 799.140 1245.300 818.220 1246.900 ;
        RECT 799.140 1243.500 800.740 1245.300 ;
        RECT 720.020 1241.900 800.740 1243.500 ;
        RECT 816.620 1243.500 818.220 1245.300 ;
        RECT 895.740 1245.300 913.900 1246.900 ;
        RECT 895.740 1243.500 897.340 1245.300 ;
        RECT 816.620 1241.900 897.340 1243.500 ;
        RECT 912.300 1243.500 913.900 1245.300 ;
        RECT 912.300 1241.900 1411.620 1243.500 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 31.350 1340.520 31.670 1340.580 ;
        RECT 1368.110 1340.520 1368.430 1340.580 ;
        RECT 31.350 1340.380 1368.430 1340.520 ;
        RECT 31.350 1340.320 31.670 1340.380 ;
        RECT 1368.110 1340.320 1368.430 1340.380 ;
        RECT 16.630 827.800 16.950 827.860 ;
        RECT 31.350 827.800 31.670 827.860 ;
        RECT 16.630 827.660 31.670 827.800 ;
        RECT 16.630 827.600 16.950 827.660 ;
        RECT 31.350 827.600 31.670 827.660 ;
      LAYER via ;
        RECT 31.380 1340.320 31.640 1340.580 ;
        RECT 1368.140 1340.320 1368.400 1340.580 ;
        RECT 16.660 827.600 16.920 827.860 ;
        RECT 31.380 827.600 31.640 827.860 ;
      LAYER met2 ;
        RECT 31.380 1340.290 31.640 1340.610 ;
        RECT 1368.140 1340.290 1368.400 1340.610 ;
        RECT 31.440 827.890 31.580 1340.290 ;
        RECT 1368.200 1325.025 1368.340 1340.290 ;
        RECT 1368.090 1321.025 1368.370 1325.025 ;
        RECT 16.660 827.570 16.920 827.890 ;
        RECT 31.380 827.570 31.640 827.890 ;
        RECT 16.720 825.365 16.860 827.570 ;
        RECT 16.650 824.995 16.930 825.365 ;
      LAYER via2 ;
        RECT 16.650 825.040 16.930 825.320 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 16.625 825.330 16.955 825.345 ;
        RECT -4.800 825.030 16.955 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 16.625 825.015 16.955 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.890 752.320 31.210 752.380 ;
        RECT 296.770 752.320 297.090 752.380 ;
        RECT 30.890 752.180 297.090 752.320 ;
        RECT 30.890 752.120 31.210 752.180 ;
        RECT 296.770 752.120 297.090 752.180 ;
        RECT 13.870 610.880 14.190 610.940 ;
        RECT 30.890 610.880 31.210 610.940 ;
        RECT 13.870 610.740 31.210 610.880 ;
        RECT 13.870 610.680 14.190 610.740 ;
        RECT 30.890 610.680 31.210 610.740 ;
      LAYER via ;
        RECT 30.920 752.120 31.180 752.380 ;
        RECT 296.800 752.120 297.060 752.380 ;
        RECT 13.900 610.680 14.160 610.940 ;
        RECT 30.920 610.680 31.180 610.940 ;
      LAYER met2 ;
        RECT 296.790 753.595 297.070 753.965 ;
        RECT 296.860 752.410 297.000 753.595 ;
        RECT 30.920 752.090 31.180 752.410 ;
        RECT 296.800 752.090 297.060 752.410 ;
        RECT 30.980 610.970 31.120 752.090 ;
        RECT 13.900 610.650 14.160 610.970 ;
        RECT 30.920 610.650 31.180 610.970 ;
        RECT 13.960 610.485 14.100 610.650 ;
        RECT 13.890 610.115 14.170 610.485 ;
      LAYER via2 ;
        RECT 296.790 753.640 297.070 753.920 ;
        RECT 13.890 610.160 14.170 610.440 ;
      LAYER met3 ;
        RECT 296.765 753.930 297.095 753.945 ;
        RECT 296.765 753.840 310.500 753.930 ;
        RECT 296.765 753.630 314.000 753.840 ;
        RECT 296.765 753.615 297.095 753.630 ;
        RECT 310.000 753.240 314.000 753.630 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 13.865 610.450 14.195 610.465 ;
        RECT -4.800 610.150 14.195 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 13.865 610.135 14.195 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 279.290 1341.200 279.610 1341.260 ;
        RECT 1071.870 1341.200 1072.190 1341.260 ;
        RECT 279.290 1341.060 1072.190 1341.200 ;
        RECT 279.290 1341.000 279.610 1341.060 ;
        RECT 1071.870 1341.000 1072.190 1341.060 ;
        RECT 19.850 400.080 20.170 400.140 ;
        RECT 279.290 400.080 279.610 400.140 ;
        RECT 19.850 399.940 279.610 400.080 ;
        RECT 19.850 399.880 20.170 399.940 ;
        RECT 279.290 399.880 279.610 399.940 ;
      LAYER via ;
        RECT 279.320 1341.000 279.580 1341.260 ;
        RECT 1071.900 1341.000 1072.160 1341.260 ;
        RECT 19.880 399.880 20.140 400.140 ;
        RECT 279.320 399.880 279.580 400.140 ;
      LAYER met2 ;
        RECT 279.320 1340.970 279.580 1341.290 ;
        RECT 1071.900 1340.970 1072.160 1341.290 ;
        RECT 279.380 400.170 279.520 1340.970 ;
        RECT 1071.960 1325.025 1072.100 1340.970 ;
        RECT 1071.850 1321.025 1072.130 1325.025 ;
        RECT 19.880 399.850 20.140 400.170 ;
        RECT 279.320 399.850 279.580 400.170 ;
        RECT 19.940 394.925 20.080 399.850 ;
        RECT 19.870 394.555 20.150 394.925 ;
      LAYER via2 ;
        RECT 19.870 394.600 20.150 394.880 ;
      LAYER met3 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 19.845 394.890 20.175 394.905 ;
        RECT -4.800 394.590 20.175 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 19.845 394.575 20.175 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1418.250 407.220 1418.570 407.280 ;
        RECT 1432.510 407.220 1432.830 407.280 ;
        RECT 1418.250 407.080 1432.830 407.220 ;
        RECT 1418.250 407.020 1418.570 407.080 ;
        RECT 1432.510 407.020 1432.830 407.080 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 1432.510 179.420 1432.830 179.480 ;
        RECT 17.090 179.280 1432.830 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 1432.510 179.220 1432.830 179.280 ;
      LAYER via ;
        RECT 1418.280 407.020 1418.540 407.280 ;
        RECT 1432.540 407.020 1432.800 407.280 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 1432.540 179.220 1432.800 179.480 ;
      LAYER met2 ;
        RECT 1418.270 409.515 1418.550 409.885 ;
        RECT 1418.340 407.310 1418.480 409.515 ;
        RECT 1418.280 406.990 1418.540 407.310 ;
        RECT 1432.540 406.990 1432.800 407.310 ;
        RECT 1432.600 179.510 1432.740 406.990 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 1432.540 179.190 1432.800 179.510 ;
      LAYER via2 ;
        RECT 1418.270 409.560 1418.550 409.840 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 1418.245 409.850 1418.575 409.865 ;
        RECT 1408.060 409.760 1418.575 409.850 ;
        RECT 1404.305 409.550 1418.575 409.760 ;
        RECT 1404.305 409.160 1408.305 409.550 ;
        RECT 1418.245 409.535 1418.575 409.550 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2114.690 787.000 2115.010 787.060 ;
        RECT 2899.450 787.000 2899.770 787.060 ;
        RECT 2114.690 786.860 2899.770 787.000 ;
        RECT 2114.690 786.800 2115.010 786.860 ;
        RECT 2899.450 786.800 2899.770 786.860 ;
        RECT 1419.170 724.440 1419.490 724.500 ;
        RECT 2114.690 724.440 2115.010 724.500 ;
        RECT 1419.170 724.300 2115.010 724.440 ;
        RECT 1419.170 724.240 1419.490 724.300 ;
        RECT 2114.690 724.240 2115.010 724.300 ;
      LAYER via ;
        RECT 2114.720 786.800 2114.980 787.060 ;
        RECT 2899.480 786.800 2899.740 787.060 ;
        RECT 1419.200 724.240 1419.460 724.500 ;
        RECT 2114.720 724.240 2114.980 724.500 ;
      LAYER met2 ;
        RECT 2899.470 791.675 2899.750 792.045 ;
        RECT 2899.540 787.090 2899.680 791.675 ;
        RECT 2114.720 786.770 2114.980 787.090 ;
        RECT 2899.480 786.770 2899.740 787.090 ;
        RECT 2114.780 724.530 2114.920 786.770 ;
        RECT 1419.200 724.210 1419.460 724.530 ;
        RECT 2114.720 724.210 2114.980 724.530 ;
        RECT 1419.260 724.045 1419.400 724.210 ;
        RECT 1419.190 723.675 1419.470 724.045 ;
      LAYER via2 ;
        RECT 2899.470 791.720 2899.750 792.000 ;
        RECT 1419.190 723.720 1419.470 724.000 ;
      LAYER met3 ;
        RECT 2899.445 792.010 2899.775 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2899.445 791.710 2924.800 792.010 ;
        RECT 2899.445 791.695 2899.775 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 1419.165 724.010 1419.495 724.025 ;
        RECT 1408.060 723.920 1419.495 724.010 ;
        RECT 1404.305 723.710 1419.495 723.920 ;
        RECT 1404.305 723.320 1408.305 723.710 ;
        RECT 1419.165 723.695 1419.495 723.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1521.750 1021.600 1522.070 1021.660 ;
        RECT 2899.450 1021.600 2899.770 1021.660 ;
        RECT 1521.750 1021.460 2899.770 1021.600 ;
        RECT 1521.750 1021.400 1522.070 1021.460 ;
        RECT 2899.450 1021.400 2899.770 1021.460 ;
        RECT 1419.170 310.320 1419.490 310.380 ;
        RECT 1521.750 310.320 1522.070 310.380 ;
        RECT 1419.170 310.180 1522.070 310.320 ;
        RECT 1419.170 310.120 1419.490 310.180 ;
        RECT 1521.750 310.120 1522.070 310.180 ;
      LAYER via ;
        RECT 1521.780 1021.400 1522.040 1021.660 ;
        RECT 2899.480 1021.400 2899.740 1021.660 ;
        RECT 1419.200 310.120 1419.460 310.380 ;
        RECT 1521.780 310.120 1522.040 310.380 ;
      LAYER met2 ;
        RECT 2899.470 1026.275 2899.750 1026.645 ;
        RECT 2899.540 1021.690 2899.680 1026.275 ;
        RECT 1521.780 1021.370 1522.040 1021.690 ;
        RECT 2899.480 1021.370 2899.740 1021.690 ;
        RECT 1521.840 310.410 1521.980 1021.370 ;
        RECT 1419.200 310.090 1419.460 310.410 ;
        RECT 1521.780 310.090 1522.040 310.410 ;
        RECT 1419.260 307.885 1419.400 310.090 ;
        RECT 1419.190 307.515 1419.470 307.885 ;
      LAYER via2 ;
        RECT 2899.470 1026.320 2899.750 1026.600 ;
        RECT 1419.190 307.560 1419.470 307.840 ;
      LAYER met3 ;
        RECT 2899.445 1026.610 2899.775 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2899.445 1026.310 2924.800 1026.610 ;
        RECT 2899.445 1026.295 2899.775 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 1419.165 307.850 1419.495 307.865 ;
        RECT 1408.060 307.760 1419.495 307.850 ;
        RECT 1404.305 307.550 1419.495 307.760 ;
        RECT 1404.305 307.160 1408.305 307.550 ;
        RECT 1419.165 307.535 1419.495 307.550 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 301.370 1314.000 301.690 1314.060 ;
        RECT 1432.970 1314.000 1433.290 1314.060 ;
        RECT 301.370 1313.860 1433.290 1314.000 ;
        RECT 301.370 1313.800 301.690 1313.860 ;
        RECT 1432.970 1313.800 1433.290 1313.860 ;
        RECT 1432.970 1262.660 1433.290 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 1432.970 1262.520 2899.310 1262.660 ;
        RECT 1432.970 1262.460 1433.290 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 301.400 1313.800 301.660 1314.060 ;
        RECT 1433.000 1313.800 1433.260 1314.060 ;
        RECT 1433.000 1262.460 1433.260 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 301.400 1313.770 301.660 1314.090 ;
        RECT 1433.000 1313.770 1433.260 1314.090 ;
        RECT 301.460 951.165 301.600 1313.770 ;
        RECT 1433.060 1262.750 1433.200 1313.770 ;
        RECT 1433.000 1262.430 1433.260 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
        RECT 301.390 950.795 301.670 951.165 ;
      LAYER via2 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
        RECT 301.390 950.840 301.670 951.120 ;
      LAYER met3 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 301.365 951.130 301.695 951.145 ;
        RECT 301.365 951.040 310.500 951.130 ;
        RECT 301.365 950.830 314.000 951.040 ;
        RECT 301.365 950.815 301.695 950.830 ;
        RECT 310.000 950.440 314.000 950.830 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1082.910 1490.800 1083.230 1490.860 ;
        RECT 2900.830 1490.800 2901.150 1490.860 ;
        RECT 1082.910 1490.660 2901.150 1490.800 ;
        RECT 1082.910 1490.600 1083.230 1490.660 ;
        RECT 2900.830 1490.600 2901.150 1490.660 ;
      LAYER via ;
        RECT 1082.940 1490.600 1083.200 1490.860 ;
        RECT 2900.860 1490.600 2901.120 1490.860 ;
      LAYER met2 ;
        RECT 2900.850 1495.475 2901.130 1495.845 ;
        RECT 2900.920 1490.890 2901.060 1495.475 ;
        RECT 1082.940 1490.570 1083.200 1490.890 ;
        RECT 2900.860 1490.570 2901.120 1490.890 ;
        RECT 1083.000 1325.050 1083.140 1490.570 ;
        RECT 1081.230 1325.025 1083.140 1325.050 ;
        RECT 1081.050 1324.910 1083.140 1325.025 ;
        RECT 1081.050 1321.025 1081.330 1324.910 ;
      LAYER via2 ;
        RECT 2900.850 1495.520 2901.130 1495.800 ;
      LAYER met3 ;
        RECT 2900.825 1495.810 2901.155 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2900.825 1495.510 2924.800 1495.810 ;
        RECT 2900.825 1495.495 2901.155 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1425.610 1725.400 1425.930 1725.460 ;
        RECT 2900.830 1725.400 2901.150 1725.460 ;
        RECT 1425.610 1725.260 2901.150 1725.400 ;
        RECT 1425.610 1725.200 1425.930 1725.260 ;
        RECT 2900.830 1725.200 2901.150 1725.260 ;
        RECT 471.110 213.420 471.430 213.480 ;
        RECT 1425.610 213.420 1425.930 213.480 ;
        RECT 471.110 213.280 1425.930 213.420 ;
        RECT 471.110 213.220 471.430 213.280 ;
        RECT 1425.610 213.220 1425.930 213.280 ;
      LAYER via ;
        RECT 1425.640 1725.200 1425.900 1725.460 ;
        RECT 2900.860 1725.200 2901.120 1725.460 ;
        RECT 471.140 213.220 471.400 213.480 ;
        RECT 1425.640 213.220 1425.900 213.480 ;
      LAYER met2 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
        RECT 2900.920 1725.490 2901.060 1730.075 ;
        RECT 1425.640 1725.170 1425.900 1725.490 ;
        RECT 2900.860 1725.170 2901.120 1725.490 ;
        RECT 471.090 216.000 471.370 220.000 ;
        RECT 471.200 213.510 471.340 216.000 ;
        RECT 1425.700 213.510 1425.840 1725.170 ;
        RECT 471.140 213.190 471.400 213.510 ;
        RECT 1425.640 213.190 1425.900 213.510 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
      LAYER met3 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1432.050 1960.000 1432.370 1960.060 ;
        RECT 2900.830 1960.000 2901.150 1960.060 ;
        RECT 1432.050 1959.860 2901.150 1960.000 ;
        RECT 1432.050 1959.800 1432.370 1959.860 ;
        RECT 2900.830 1959.800 2901.150 1959.860 ;
        RECT 1242.070 213.760 1242.390 213.820 ;
        RECT 1432.050 213.760 1432.370 213.820 ;
        RECT 1242.070 213.620 1432.370 213.760 ;
        RECT 1242.070 213.560 1242.390 213.620 ;
        RECT 1432.050 213.560 1432.370 213.620 ;
      LAYER via ;
        RECT 1432.080 1959.800 1432.340 1960.060 ;
        RECT 2900.860 1959.800 2901.120 1960.060 ;
        RECT 1242.100 213.560 1242.360 213.820 ;
        RECT 1432.080 213.560 1432.340 213.820 ;
      LAYER met2 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
        RECT 2900.920 1960.090 2901.060 1964.675 ;
        RECT 1432.080 1959.770 1432.340 1960.090 ;
        RECT 2900.860 1959.770 2901.120 1960.090 ;
        RECT 1242.050 216.000 1242.330 220.000 ;
        RECT 1242.160 213.850 1242.300 216.000 ;
        RECT 1432.140 213.850 1432.280 1959.770 ;
        RECT 1242.100 213.530 1242.360 213.850 ;
        RECT 1432.080 213.530 1432.340 213.850 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
      LAYER met3 ;
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 312.410 2194.600 312.730 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 312.410 2194.460 2901.150 2194.600 ;
        RECT 312.410 2194.400 312.730 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
        RECT 303.210 641.820 303.530 641.880 ;
        RECT 311.950 641.820 312.270 641.880 ;
        RECT 303.210 641.680 312.270 641.820 ;
        RECT 303.210 641.620 303.530 641.680 ;
        RECT 311.950 641.620 312.270 641.680 ;
      LAYER via ;
        RECT 312.440 2194.400 312.700 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
        RECT 303.240 641.620 303.500 641.880 ;
        RECT 311.980 641.620 312.240 641.880 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 312.440 2194.370 312.700 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 303.240 641.590 303.500 641.910 ;
        RECT 311.980 641.820 312.240 641.910 ;
        RECT 312.500 641.820 312.640 2194.370 ;
        RECT 311.980 641.680 312.640 641.820 ;
        RECT 311.980 641.590 312.240 641.680 ;
        RECT 303.300 556.765 303.440 641.590 ;
        RECT 303.230 556.395 303.510 556.765 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 303.230 556.440 303.510 556.720 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 303.205 556.730 303.535 556.745 ;
        RECT 303.205 556.640 310.500 556.730 ;
        RECT 303.205 556.430 314.000 556.640 ;
        RECT 303.205 556.415 303.535 556.430 ;
        RECT 310.000 556.040 314.000 556.430 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 289.920 1419.490 289.980 ;
        RECT 2473.490 289.920 2473.810 289.980 ;
        RECT 1419.170 289.780 2473.810 289.920 ;
        RECT 1419.170 289.720 1419.490 289.780 ;
        RECT 2473.490 289.720 2473.810 289.780 ;
        RECT 2473.490 206.960 2473.810 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2473.490 206.820 2901.150 206.960 ;
        RECT 2473.490 206.760 2473.810 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 1419.200 289.720 1419.460 289.980 ;
        RECT 2473.520 289.720 2473.780 289.980 ;
        RECT 2473.520 206.760 2473.780 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 1419.190 292.555 1419.470 292.925 ;
        RECT 1419.260 290.010 1419.400 292.555 ;
        RECT 1419.200 289.690 1419.460 290.010 ;
        RECT 2473.520 289.690 2473.780 290.010 ;
        RECT 2473.580 207.050 2473.720 289.690 ;
        RECT 2473.520 206.730 2473.780 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 1419.190 292.600 1419.470 292.880 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 1419.165 292.890 1419.495 292.905 ;
        RECT 1408.060 292.800 1419.495 292.890 ;
        RECT 1404.305 292.590 1419.495 292.800 ;
        RECT 1404.305 292.200 1408.305 292.590 ;
        RECT 1419.165 292.575 1419.495 292.590 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1425.150 2546.500 1425.470 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 1425.150 2546.360 2901.150 2546.500 ;
        RECT 1425.150 2546.300 1425.470 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
      LAYER via ;
        RECT 1425.180 2546.300 1425.440 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 1425.180 2546.270 1425.440 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 950.410 216.000 950.690 220.000 ;
        RECT 950.520 209.965 950.660 216.000 ;
        RECT 1425.240 209.965 1425.380 2546.270 ;
        RECT 950.450 209.595 950.730 209.965 ;
        RECT 1425.170 209.595 1425.450 209.965 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
        RECT 950.450 209.640 950.730 209.920 ;
        RECT 1425.170 209.640 1425.450 209.920 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 950.425 209.930 950.755 209.945 ;
        RECT 1425.145 209.930 1425.475 209.945 ;
        RECT 950.425 209.630 1425.475 209.930 ;
        RECT 950.425 209.615 950.755 209.630 ;
        RECT 1425.145 209.615 1425.475 209.630 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2608.270 2782.120 2608.590 2782.180 ;
        RECT 2646.450 2782.120 2646.770 2782.180 ;
        RECT 2608.270 2781.980 2646.770 2782.120 ;
        RECT 2608.270 2781.920 2608.590 2781.980 ;
        RECT 2646.450 2781.920 2646.770 2781.980 ;
        RECT 2076.970 2781.780 2077.290 2781.840 ;
        RECT 2124.350 2781.780 2124.670 2781.840 ;
        RECT 2076.970 2781.640 2124.670 2781.780 ;
        RECT 2076.970 2781.580 2077.290 2781.640 ;
        RECT 2124.350 2781.580 2124.670 2781.640 ;
      LAYER via ;
        RECT 2608.300 2781.920 2608.560 2782.180 ;
        RECT 2646.480 2781.920 2646.740 2782.180 ;
        RECT 2077.000 2781.580 2077.260 2781.840 ;
        RECT 2124.380 2781.580 2124.640 2781.840 ;
      LAYER met2 ;
        RECT 2670.390 2782.715 2670.670 2783.085 ;
        RECT 2704.890 2782.715 2705.170 2783.085 ;
        RECT 2124.370 2782.035 2124.650 2782.405 ;
        RECT 2125.290 2782.035 2125.570 2782.405 ;
        RECT 2608.290 2782.035 2608.570 2782.405 ;
        RECT 2124.440 2781.870 2124.580 2782.035 ;
        RECT 2077.000 2781.725 2077.260 2781.870 ;
        RECT 2076.990 2781.355 2077.270 2781.725 ;
        RECT 2124.380 2781.550 2124.640 2781.870 ;
        RECT 2125.360 2779.685 2125.500 2782.035 ;
        RECT 2608.300 2781.890 2608.560 2782.035 ;
        RECT 2646.480 2781.890 2646.740 2782.210 ;
        RECT 2646.540 2781.045 2646.680 2781.890 ;
        RECT 2646.470 2780.675 2646.750 2781.045 ;
        RECT 2669.930 2780.930 2670.210 2781.045 ;
        RECT 2670.460 2780.930 2670.600 2782.715 ;
        RECT 2704.960 2781.045 2705.100 2782.715 ;
        RECT 2766.990 2782.290 2767.270 2782.405 ;
        RECT 2766.600 2782.150 2767.270 2782.290 ;
        RECT 2766.600 2781.725 2766.740 2782.150 ;
        RECT 2766.990 2782.035 2767.270 2782.150 ;
        RECT 2766.530 2781.355 2766.810 2781.725 ;
        RECT 2669.930 2780.790 2670.600 2780.930 ;
        RECT 2669.930 2780.675 2670.210 2780.790 ;
        RECT 2704.890 2780.675 2705.170 2781.045 ;
        RECT 2125.290 2779.315 2125.570 2779.685 ;
        RECT 431.530 216.000 431.810 220.000 ;
        RECT 431.640 213.365 431.780 216.000 ;
        RECT 431.570 212.995 431.850 213.365 ;
      LAYER via2 ;
        RECT 2670.390 2782.760 2670.670 2783.040 ;
        RECT 2704.890 2782.760 2705.170 2783.040 ;
        RECT 2124.370 2782.080 2124.650 2782.360 ;
        RECT 2125.290 2782.080 2125.570 2782.360 ;
        RECT 2608.290 2782.080 2608.570 2782.360 ;
        RECT 2076.990 2781.400 2077.270 2781.680 ;
        RECT 2646.470 2780.720 2646.750 2781.000 ;
        RECT 2669.930 2780.720 2670.210 2781.000 ;
        RECT 2766.990 2782.080 2767.270 2782.360 ;
        RECT 2766.530 2781.400 2766.810 2781.680 ;
        RECT 2704.890 2780.720 2705.170 2781.000 ;
        RECT 2125.290 2779.360 2125.570 2779.640 ;
        RECT 431.570 213.040 431.850 213.320 ;
      LAYER met3 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2916.710 2786.150 2924.800 2786.450 ;
        RECT 2670.365 2783.050 2670.695 2783.065 ;
        RECT 2704.865 2783.050 2705.195 2783.065 ;
        RECT 2670.365 2782.750 2705.195 2783.050 ;
        RECT 2670.365 2782.735 2670.695 2782.750 ;
        RECT 2704.865 2782.735 2705.195 2782.750 ;
        RECT 1497.110 2782.370 1497.490 2782.380 ;
        RECT 2124.345 2782.370 2124.675 2782.385 ;
        RECT 2125.265 2782.370 2125.595 2782.385 ;
        RECT 1435.510 2782.070 1463.410 2782.370 ;
        RECT 1430.870 2781.010 1431.250 2781.020 ;
        RECT 1435.510 2781.010 1435.810 2782.070 ;
        RECT 1430.870 2780.710 1435.810 2781.010 ;
        RECT 1463.110 2781.010 1463.410 2782.070 ;
        RECT 1497.110 2782.070 1580.250 2782.370 ;
        RECT 1497.110 2782.060 1497.490 2782.070 ;
        RECT 1579.950 2781.690 1580.250 2782.070 ;
        RECT 1628.710 2782.070 1676.850 2782.370 ;
        RECT 1579.950 2781.390 1628.090 2781.690 ;
        RECT 1497.110 2781.010 1497.490 2781.020 ;
        RECT 1463.110 2780.710 1497.490 2781.010 ;
        RECT 1627.790 2781.010 1628.090 2781.390 ;
        RECT 1628.710 2781.010 1629.010 2782.070 ;
        RECT 1676.550 2781.690 1676.850 2782.070 ;
        RECT 1725.310 2782.070 1773.450 2782.370 ;
        RECT 1676.550 2781.390 1724.690 2781.690 ;
        RECT 1627.790 2780.710 1629.010 2781.010 ;
        RECT 1724.390 2781.010 1724.690 2781.390 ;
        RECT 1725.310 2781.010 1725.610 2782.070 ;
        RECT 1773.150 2781.690 1773.450 2782.070 ;
        RECT 1821.910 2782.070 1870.050 2782.370 ;
        RECT 1773.150 2781.390 1821.290 2781.690 ;
        RECT 1724.390 2780.710 1725.610 2781.010 ;
        RECT 1820.990 2781.010 1821.290 2781.390 ;
        RECT 1821.910 2781.010 1822.210 2782.070 ;
        RECT 1869.750 2781.690 1870.050 2782.070 ;
        RECT 1918.510 2782.070 1966.650 2782.370 ;
        RECT 1869.750 2781.390 1917.890 2781.690 ;
        RECT 1820.990 2780.710 1822.210 2781.010 ;
        RECT 1917.590 2781.010 1917.890 2781.390 ;
        RECT 1918.510 2781.010 1918.810 2782.070 ;
        RECT 1966.350 2781.690 1966.650 2782.070 ;
        RECT 2015.110 2782.070 2063.250 2782.370 ;
        RECT 1966.350 2781.390 2014.490 2781.690 ;
        RECT 1917.590 2780.710 1918.810 2781.010 ;
        RECT 2014.190 2781.010 2014.490 2781.390 ;
        RECT 2015.110 2781.010 2015.410 2782.070 ;
        RECT 2062.950 2781.690 2063.250 2782.070 ;
        RECT 2124.345 2782.070 2125.595 2782.370 ;
        RECT 2124.345 2782.055 2124.675 2782.070 ;
        RECT 2125.265 2782.055 2125.595 2782.070 ;
        RECT 2173.310 2782.370 2173.690 2782.380 ;
        RECT 2608.265 2782.370 2608.595 2782.385 ;
        RECT 2173.310 2782.070 2256.450 2782.370 ;
        RECT 2173.310 2782.060 2173.690 2782.070 ;
        RECT 2076.965 2781.690 2077.295 2781.705 ;
        RECT 2062.950 2781.390 2077.295 2781.690 ;
        RECT 2256.150 2781.690 2256.450 2782.070 ;
        RECT 2304.910 2782.070 2353.050 2782.370 ;
        RECT 2256.150 2781.390 2304.290 2781.690 ;
        RECT 2076.965 2781.375 2077.295 2781.390 ;
        RECT 2014.190 2780.710 2015.410 2781.010 ;
        RECT 2303.990 2781.010 2304.290 2781.390 ;
        RECT 2304.910 2781.010 2305.210 2782.070 ;
        RECT 2352.750 2781.690 2353.050 2782.070 ;
        RECT 2401.510 2782.070 2449.650 2782.370 ;
        RECT 2352.750 2781.390 2400.890 2781.690 ;
        RECT 2303.990 2780.710 2305.210 2781.010 ;
        RECT 2400.590 2781.010 2400.890 2781.390 ;
        RECT 2401.510 2781.010 2401.810 2782.070 ;
        RECT 2449.350 2781.690 2449.650 2782.070 ;
        RECT 2498.110 2782.070 2546.250 2782.370 ;
        RECT 2449.350 2781.390 2497.490 2781.690 ;
        RECT 2400.590 2780.710 2401.810 2781.010 ;
        RECT 2497.190 2781.010 2497.490 2781.390 ;
        RECT 2498.110 2781.010 2498.410 2782.070 ;
        RECT 2545.950 2781.690 2546.250 2782.070 ;
        RECT 2594.710 2782.070 2608.595 2782.370 ;
        RECT 2545.950 2781.390 2594.090 2781.690 ;
        RECT 2497.190 2780.710 2498.410 2781.010 ;
        RECT 2593.790 2781.010 2594.090 2781.390 ;
        RECT 2594.710 2781.010 2595.010 2782.070 ;
        RECT 2608.265 2782.055 2608.595 2782.070 ;
        RECT 2766.965 2782.370 2767.295 2782.385 ;
        RECT 2766.965 2782.070 2836.050 2782.370 ;
        RECT 2766.965 2782.055 2767.295 2782.070 ;
        RECT 2766.505 2781.690 2766.835 2781.705 ;
        RECT 2752.950 2781.390 2766.835 2781.690 ;
        RECT 2835.750 2781.690 2836.050 2782.070 ;
        RECT 2916.710 2781.690 2917.010 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2835.750 2781.390 2883.890 2781.690 ;
        RECT 2593.790 2780.710 2595.010 2781.010 ;
        RECT 2646.445 2781.010 2646.775 2781.025 ;
        RECT 2669.905 2781.010 2670.235 2781.025 ;
        RECT 2646.445 2780.710 2670.235 2781.010 ;
        RECT 1430.870 2780.700 1431.250 2780.710 ;
        RECT 1497.110 2780.700 1497.490 2780.710 ;
        RECT 2646.445 2780.695 2646.775 2780.710 ;
        RECT 2669.905 2780.695 2670.235 2780.710 ;
        RECT 2704.865 2781.010 2705.195 2781.025 ;
        RECT 2752.950 2781.010 2753.250 2781.390 ;
        RECT 2766.505 2781.375 2766.835 2781.390 ;
        RECT 2704.865 2780.710 2753.250 2781.010 ;
        RECT 2883.590 2781.010 2883.890 2781.390 ;
        RECT 2884.510 2781.390 2917.010 2781.690 ;
        RECT 2884.510 2781.010 2884.810 2781.390 ;
        RECT 2883.590 2780.710 2884.810 2781.010 ;
        RECT 2704.865 2780.695 2705.195 2780.710 ;
        RECT 2125.265 2779.650 2125.595 2779.665 ;
        RECT 2173.310 2779.650 2173.690 2779.660 ;
        RECT 2125.265 2779.350 2173.690 2779.650 ;
        RECT 2125.265 2779.335 2125.595 2779.350 ;
        RECT 2173.310 2779.340 2173.690 2779.350 ;
        RECT 431.545 213.330 431.875 213.345 ;
        RECT 1430.870 213.330 1431.250 213.340 ;
        RECT 431.545 213.030 1431.250 213.330 ;
        RECT 431.545 213.015 431.875 213.030 ;
        RECT 1430.870 213.020 1431.250 213.030 ;
      LAYER via3 ;
        RECT 1430.900 2780.700 1431.220 2781.020 ;
        RECT 1497.140 2782.060 1497.460 2782.380 ;
        RECT 1497.140 2780.700 1497.460 2781.020 ;
        RECT 2173.340 2782.060 2173.660 2782.380 ;
        RECT 2173.340 2779.340 2173.660 2779.660 ;
        RECT 1430.900 213.020 1431.220 213.340 ;
      LAYER met4 ;
        RECT 1497.135 2782.055 1497.465 2782.385 ;
        RECT 2173.335 2782.055 2173.665 2782.385 ;
        RECT 1497.150 2781.025 1497.450 2782.055 ;
        RECT 1430.895 2780.695 1431.225 2781.025 ;
        RECT 1497.135 2780.695 1497.465 2781.025 ;
        RECT 1430.910 213.345 1431.210 2780.695 ;
        RECT 2173.350 2779.665 2173.650 2782.055 ;
        RECT 2173.335 2779.335 2173.665 2779.665 ;
        RECT 1430.895 213.015 1431.225 213.345 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1117.410 3015.700 1117.730 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 1117.410 3015.560 2901.150 3015.700 ;
        RECT 1117.410 3015.500 1117.730 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 1117.440 3015.500 1117.700 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 1117.440 3015.470 1117.700 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 1117.500 1325.050 1117.640 3015.470 ;
        RECT 1116.190 1325.025 1117.640 1325.050 ;
        RECT 1116.010 1324.910 1117.640 1325.025 ;
        RECT 1116.010 1321.025 1116.290 1324.910 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1569.590 3250.300 1569.910 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1569.590 3250.160 2901.150 3250.300 ;
        RECT 1569.590 3250.100 1569.910 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 1421.010 710.500 1421.330 710.560 ;
        RECT 1569.590 710.500 1569.910 710.560 ;
        RECT 1421.010 710.360 1569.910 710.500 ;
        RECT 1421.010 710.300 1421.330 710.360 ;
        RECT 1569.590 710.300 1569.910 710.360 ;
      LAYER via ;
        RECT 1569.620 3250.100 1569.880 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 1421.040 710.300 1421.300 710.560 ;
        RECT 1569.620 710.300 1569.880 710.560 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1569.620 3250.070 1569.880 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1569.680 710.590 1569.820 3250.070 ;
        RECT 1421.040 710.445 1421.300 710.590 ;
        RECT 1421.030 710.075 1421.310 710.445 ;
        RECT 1569.620 710.270 1569.880 710.590 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
        RECT 1421.030 710.120 1421.310 710.400 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 1421.005 710.410 1421.335 710.425 ;
        RECT 1408.060 710.320 1421.335 710.410 ;
        RECT 1404.305 710.110 1421.335 710.320 ;
        RECT 1404.305 709.720 1408.305 710.110 ;
        RECT 1421.005 710.095 1421.335 710.110 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1597.190 3484.900 1597.510 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1597.190 3484.760 2901.150 3484.900 ;
        RECT 1597.190 3484.700 1597.510 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 1419.170 1193.640 1419.490 1193.700 ;
        RECT 1597.190 1193.640 1597.510 1193.700 ;
        RECT 1419.170 1193.500 1597.510 1193.640 ;
        RECT 1419.170 1193.440 1419.490 1193.500 ;
        RECT 1597.190 1193.440 1597.510 1193.500 ;
      LAYER via ;
        RECT 1597.220 3484.700 1597.480 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 1419.200 1193.440 1419.460 1193.700 ;
        RECT 1597.220 1193.440 1597.480 1193.700 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1597.220 3484.670 1597.480 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1597.280 1193.730 1597.420 3484.670 ;
        RECT 1419.200 1193.410 1419.460 1193.730 ;
        RECT 1597.220 1193.410 1597.480 1193.730 ;
        RECT 1419.260 1191.885 1419.400 1193.410 ;
        RECT 1419.190 1191.515 1419.470 1191.885 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 1419.190 1191.560 1419.470 1191.840 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 1419.165 1191.850 1419.495 1191.865 ;
        RECT 1408.060 1191.760 1419.495 1191.850 ;
        RECT 1404.305 1191.550 1419.495 1191.760 ;
        RECT 1404.305 1191.160 1408.305 1191.550 ;
        RECT 1419.165 1191.535 1419.495 1191.550 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.590 1355.820 304.910 1355.880 ;
        RECT 2635.870 1355.820 2636.190 1355.880 ;
        RECT 304.590 1355.680 2636.190 1355.820 ;
        RECT 304.590 1355.620 304.910 1355.680 ;
        RECT 2635.870 1355.620 2636.190 1355.680 ;
      LAYER via ;
        RECT 304.620 1355.620 304.880 1355.880 ;
        RECT 2635.900 1355.620 2636.160 1355.880 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 1355.910 2636.100 3517.600 ;
        RECT 304.620 1355.590 304.880 1355.910 ;
        RECT 2635.900 1355.590 2636.160 1355.910 ;
        RECT 304.680 1191.885 304.820 1355.590 ;
        RECT 304.610 1191.515 304.890 1191.885 ;
      LAYER via2 ;
        RECT 304.610 1191.560 304.890 1191.840 ;
      LAYER met3 ;
        RECT 304.585 1191.850 304.915 1191.865 ;
        RECT 304.585 1191.760 310.500 1191.850 ;
        RECT 304.585 1191.550 314.000 1191.760 ;
        RECT 304.585 1191.535 304.915 1191.550 ;
        RECT 310.000 1191.160 314.000 1191.550 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 302.290 1362.620 302.610 1362.680 ;
        RECT 2311.570 1362.620 2311.890 1362.680 ;
        RECT 302.290 1362.480 2311.890 1362.620 ;
        RECT 302.290 1362.420 302.610 1362.480 ;
        RECT 2311.570 1362.420 2311.890 1362.480 ;
      LAYER via ;
        RECT 302.320 1362.420 302.580 1362.680 ;
        RECT 2311.600 1362.420 2311.860 1362.680 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 1362.710 2311.800 3517.600 ;
        RECT 302.320 1362.390 302.580 1362.710 ;
        RECT 2311.600 1362.390 2311.860 1362.710 ;
        RECT 302.380 1287.085 302.520 1362.390 ;
        RECT 302.310 1286.715 302.590 1287.085 ;
      LAYER via2 ;
        RECT 302.310 1286.760 302.590 1287.040 ;
      LAYER met3 ;
        RECT 302.285 1287.050 302.615 1287.065 ;
        RECT 302.285 1286.960 310.500 1287.050 ;
        RECT 302.285 1286.750 314.000 1286.960 ;
        RECT 302.285 1286.735 302.615 1286.750 ;
        RECT 310.000 1286.360 314.000 1286.750 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.010 3501.560 524.330 3501.620 ;
        RECT 1987.270 3501.560 1987.590 3501.620 ;
        RECT 524.010 3501.420 1987.590 3501.560 ;
        RECT 524.010 3501.360 524.330 3501.420 ;
        RECT 1987.270 3501.360 1987.590 3501.420 ;
      LAYER via ;
        RECT 524.040 3501.360 524.300 3501.620 ;
        RECT 1987.300 3501.360 1987.560 3501.620 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3501.650 1987.500 3517.600 ;
        RECT 524.040 3501.330 524.300 3501.650 ;
        RECT 1987.300 3501.330 1987.560 3501.650 ;
        RECT 524.100 1325.050 524.240 3501.330 ;
        RECT 522.790 1325.025 524.240 1325.050 ;
        RECT 522.610 1324.910 524.240 1325.025 ;
        RECT 522.610 1321.025 522.890 1324.910 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1438.490 3502.580 1438.810 3502.640 ;
        RECT 1662.510 3502.580 1662.830 3502.640 ;
        RECT 1438.490 3502.440 1662.830 3502.580 ;
        RECT 1438.490 3502.380 1438.810 3502.440 ;
        RECT 1662.510 3502.380 1662.830 3502.440 ;
        RECT 975.270 212.400 975.590 212.460 ;
        RECT 1438.490 212.400 1438.810 212.460 ;
        RECT 975.270 212.260 1438.810 212.400 ;
        RECT 975.270 212.200 975.590 212.260 ;
        RECT 1438.490 212.200 1438.810 212.260 ;
      LAYER via ;
        RECT 1438.520 3502.380 1438.780 3502.640 ;
        RECT 1662.540 3502.380 1662.800 3502.640 ;
        RECT 975.300 212.200 975.560 212.460 ;
        RECT 1438.520 212.200 1438.780 212.460 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3502.670 1662.740 3517.600 ;
        RECT 1438.520 3502.350 1438.780 3502.670 ;
        RECT 1662.540 3502.350 1662.800 3502.670 ;
        RECT 975.250 216.000 975.530 220.000 ;
        RECT 975.360 212.490 975.500 216.000 ;
        RECT 1438.580 212.490 1438.720 3502.350 ;
        RECT 975.300 212.170 975.560 212.490 ;
        RECT 1438.520 212.170 1438.780 212.490 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3501.845 1338.440 3517.600 ;
        RECT 1338.230 3501.475 1338.510 3501.845 ;
        RECT 841.850 216.000 842.130 220.000 ;
        RECT 841.960 205.885 842.100 216.000 ;
        RECT 841.890 205.515 842.170 205.885 ;
      LAYER via2 ;
        RECT 1338.230 3501.520 1338.510 3501.800 ;
        RECT 841.890 205.560 842.170 205.840 ;
      LAYER met3 ;
        RECT 1338.205 3501.810 1338.535 3501.825 ;
        RECT 1428.110 3501.810 1428.490 3501.820 ;
        RECT 1338.205 3501.510 1428.490 3501.810 ;
        RECT 1338.205 3501.495 1338.535 3501.510 ;
        RECT 1428.110 3501.500 1428.490 3501.510 ;
        RECT 841.865 205.850 842.195 205.865 ;
        RECT 1428.110 205.850 1428.490 205.860 ;
        RECT 841.865 205.550 1428.490 205.850 ;
        RECT 841.865 205.535 842.195 205.550 ;
        RECT 1428.110 205.540 1428.490 205.550 ;
      LAYER via3 ;
        RECT 1428.140 3501.500 1428.460 3501.820 ;
        RECT 1428.140 205.540 1428.460 205.860 ;
      LAYER met4 ;
        RECT 1428.135 3501.495 1428.465 3501.825 ;
        RECT 1428.150 205.865 1428.450 3501.495 ;
        RECT 1428.135 205.535 1428.465 205.865 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 821.340 1419.490 821.400 ;
        RECT 2507.990 821.340 2508.310 821.400 ;
        RECT 1419.170 821.200 2508.310 821.340 ;
        RECT 1419.170 821.140 1419.490 821.200 ;
        RECT 2507.990 821.140 2508.310 821.200 ;
        RECT 2507.990 441.560 2508.310 441.620 ;
        RECT 2899.450 441.560 2899.770 441.620 ;
        RECT 2507.990 441.420 2899.770 441.560 ;
        RECT 2507.990 441.360 2508.310 441.420 ;
        RECT 2899.450 441.360 2899.770 441.420 ;
      LAYER via ;
        RECT 1419.200 821.140 1419.460 821.400 ;
        RECT 2508.020 821.140 2508.280 821.400 ;
        RECT 2508.020 441.360 2508.280 441.620 ;
        RECT 2899.480 441.360 2899.740 441.620 ;
      LAYER met2 ;
        RECT 1419.190 827.035 1419.470 827.405 ;
        RECT 1419.260 821.430 1419.400 827.035 ;
        RECT 1419.200 821.110 1419.460 821.430 ;
        RECT 2508.020 821.110 2508.280 821.430 ;
        RECT 2508.080 441.650 2508.220 821.110 ;
        RECT 2508.020 441.330 2508.280 441.650 ;
        RECT 2899.480 441.330 2899.740 441.650 ;
        RECT 2899.540 439.805 2899.680 441.330 ;
        RECT 2899.470 439.435 2899.750 439.805 ;
      LAYER via2 ;
        RECT 1419.190 827.080 1419.470 827.360 ;
        RECT 2899.470 439.480 2899.750 439.760 ;
      LAYER met3 ;
        RECT 1419.165 827.370 1419.495 827.385 ;
        RECT 1408.060 827.280 1419.495 827.370 ;
        RECT 1404.305 827.070 1419.495 827.280 ;
        RECT 1404.305 826.680 1408.305 827.070 ;
        RECT 1419.165 827.055 1419.495 827.070 ;
        RECT 2899.445 439.770 2899.775 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2899.445 439.470 2924.800 439.770 ;
        RECT 2899.445 439.455 2899.775 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1013.910 1369.760 1014.230 1369.820 ;
        RECT 1417.330 1369.760 1417.650 1369.820 ;
        RECT 1013.910 1369.620 1417.650 1369.760 ;
        RECT 1013.910 1369.560 1014.230 1369.620 ;
        RECT 1417.330 1369.560 1417.650 1369.620 ;
      LAYER via ;
        RECT 1013.940 1369.560 1014.200 1369.820 ;
        RECT 1417.360 1369.560 1417.620 1369.820 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 1369.850 1014.140 3517.600 ;
        RECT 1013.940 1369.530 1014.200 1369.850 ;
        RECT 1417.360 1369.530 1417.620 1369.850 ;
        RECT 1417.420 957.965 1417.560 1369.530 ;
        RECT 1417.350 957.595 1417.630 957.965 ;
      LAYER via2 ;
        RECT 1417.350 957.640 1417.630 957.920 ;
      LAYER met3 ;
        RECT 1417.325 957.930 1417.655 957.945 ;
        RECT 1408.060 957.840 1417.655 957.930 ;
        RECT 1404.305 957.630 1417.655 957.840 ;
        RECT 1404.305 957.240 1408.305 957.630 ;
        RECT 1417.325 957.615 1417.655 957.630 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 689.150 3502.920 689.470 3502.980 ;
        RECT 1415.030 3502.920 1415.350 3502.980 ;
        RECT 689.150 3502.780 1415.350 3502.920 ;
        RECT 689.150 3502.720 689.470 3502.780 ;
        RECT 1415.030 3502.720 1415.350 3502.780 ;
      LAYER via ;
        RECT 689.180 3502.720 689.440 3502.980 ;
        RECT 1415.060 3502.720 1415.320 3502.980 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3503.010 689.380 3517.600 ;
        RECT 689.180 3502.690 689.440 3503.010 ;
        RECT 1415.060 3502.690 1415.320 3503.010 ;
        RECT 1415.120 1048.405 1415.260 3502.690 ;
        RECT 1415.050 1048.035 1415.330 1048.405 ;
        RECT 1108.650 216.000 1108.930 220.000 ;
        RECT 1108.760 205.205 1108.900 216.000 ;
        RECT 1108.690 204.835 1108.970 205.205 ;
      LAYER via2 ;
        RECT 1415.050 1048.080 1415.330 1048.360 ;
        RECT 1108.690 204.880 1108.970 205.160 ;
      LAYER met3 ;
        RECT 1415.025 1048.380 1415.355 1048.385 ;
        RECT 1415.025 1048.370 1415.610 1048.380 ;
        RECT 1414.800 1048.070 1415.610 1048.370 ;
        RECT 1415.025 1048.060 1415.610 1048.070 ;
        RECT 1415.025 1048.055 1415.355 1048.060 ;
        RECT 1108.665 205.170 1108.995 205.185 ;
        RECT 1415.230 205.170 1415.610 205.180 ;
        RECT 1108.665 204.870 1415.610 205.170 ;
        RECT 1108.665 204.855 1108.995 204.870 ;
        RECT 1415.230 204.860 1415.610 204.870 ;
      LAYER via3 ;
        RECT 1415.260 1048.060 1415.580 1048.380 ;
        RECT 1415.260 204.860 1415.580 205.180 ;
      LAYER met4 ;
        RECT 1415.255 1048.055 1415.585 1048.385 ;
        RECT 1415.270 205.185 1415.570 1048.055 ;
        RECT 1415.255 204.855 1415.585 205.185 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.580 365.170 3502.640 ;
        RECT 1345.570 3502.580 1345.890 3502.640 ;
        RECT 364.850 3502.440 1345.890 3502.580 ;
        RECT 364.850 3502.380 365.170 3502.440 ;
        RECT 1345.570 3502.380 1345.890 3502.440 ;
      LAYER via ;
        RECT 364.880 3502.380 365.140 3502.640 ;
        RECT 1345.600 3502.380 1345.860 3502.640 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3502.670 365.080 3517.600 ;
        RECT 364.880 3502.350 365.140 3502.670 ;
        RECT 1345.600 3502.350 1345.860 3502.670 ;
        RECT 1345.660 1324.370 1345.800 3502.350 ;
        RECT 1348.770 1324.370 1349.050 1325.025 ;
        RECT 1345.660 1324.230 1349.050 1324.370 ;
        RECT 1348.770 1321.025 1349.050 1324.230 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 40.625 3429.325 40.795 3477.435 ;
        RECT 40.165 2898.585 40.335 2946.355 ;
        RECT 40.165 2704.785 40.335 2752.895 ;
        RECT 40.165 1952.705 40.335 1994.695 ;
        RECT 40.165 1738.845 40.335 1786.955 ;
        RECT 40.165 1684.105 40.335 1705.015 ;
        RECT 39.705 1635.485 39.875 1683.255 ;
        RECT 40.625 1400.885 40.795 1448.995 ;
        RECT 40.165 1075.845 40.335 1110.695 ;
        RECT 39.705 965.685 39.875 1007.335 ;
        RECT 39.705 579.785 39.875 627.895 ;
        RECT 40.165 496.485 40.335 531.335 ;
      LAYER mcon ;
        RECT 40.625 3477.265 40.795 3477.435 ;
        RECT 40.165 2946.185 40.335 2946.355 ;
        RECT 40.165 2752.725 40.335 2752.895 ;
        RECT 40.165 1994.525 40.335 1994.695 ;
        RECT 40.165 1786.785 40.335 1786.955 ;
        RECT 40.165 1704.845 40.335 1705.015 ;
        RECT 39.705 1683.085 39.875 1683.255 ;
        RECT 40.625 1448.825 40.795 1448.995 ;
        RECT 40.165 1110.525 40.335 1110.695 ;
        RECT 39.705 1007.165 39.875 1007.335 ;
        RECT 39.705 627.725 39.875 627.895 ;
        RECT 40.165 531.165 40.335 531.335 ;
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 40.565 3477.420 40.855 3477.465 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 40.565 3477.280 41.330 3477.420 ;
        RECT 40.565 3477.235 40.855 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 40.355 3429.340 40.870 3429.480 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3270.700 40.410 3270.760 ;
        RECT 41.010 3270.700 41.330 3270.760 ;
        RECT 40.090 3270.560 41.330 3270.700 ;
        RECT 40.090 3270.500 40.410 3270.560 ;
        RECT 41.010 3270.500 41.330 3270.560 ;
        RECT 40.090 3174.140 40.410 3174.200 ;
        RECT 41.010 3174.140 41.330 3174.200 ;
        RECT 40.090 3174.000 41.330 3174.140 ;
        RECT 40.090 3173.940 40.410 3174.000 ;
        RECT 41.010 3173.940 41.330 3174.000 ;
        RECT 40.090 3077.580 40.410 3077.640 ;
        RECT 41.010 3077.580 41.330 3077.640 ;
        RECT 40.090 3077.440 41.330 3077.580 ;
        RECT 40.090 3077.380 40.410 3077.440 ;
        RECT 41.010 3077.380 41.330 3077.440 ;
        RECT 40.090 2981.020 40.410 2981.080 ;
        RECT 41.010 2981.020 41.330 2981.080 ;
        RECT 40.090 2980.880 41.330 2981.020 ;
        RECT 40.090 2980.820 40.410 2980.880 ;
        RECT 41.010 2980.820 41.330 2980.880 ;
        RECT 40.090 2946.340 40.410 2946.400 ;
        RECT 39.895 2946.200 40.410 2946.340 ;
        RECT 40.090 2946.140 40.410 2946.200 ;
        RECT 40.090 2898.740 40.410 2898.800 ;
        RECT 39.895 2898.600 40.410 2898.740 ;
        RECT 40.090 2898.540 40.410 2898.600 ;
        RECT 39.630 2898.060 39.950 2898.120 ;
        RECT 40.550 2898.060 40.870 2898.120 ;
        RECT 39.630 2897.920 40.870 2898.060 ;
        RECT 39.630 2897.860 39.950 2897.920 ;
        RECT 40.550 2897.860 40.870 2897.920 ;
        RECT 39.630 2814.760 39.950 2814.820 ;
        RECT 40.550 2814.760 40.870 2814.820 ;
        RECT 39.630 2814.620 40.870 2814.760 ;
        RECT 39.630 2814.560 39.950 2814.620 ;
        RECT 40.550 2814.560 40.870 2814.620 ;
        RECT 40.090 2752.880 40.410 2752.940 ;
        RECT 39.895 2752.740 40.410 2752.880 ;
        RECT 40.090 2752.680 40.410 2752.740 ;
        RECT 40.105 2704.940 40.395 2704.985 ;
        RECT 41.010 2704.940 41.330 2705.000 ;
        RECT 40.105 2704.800 41.330 2704.940 ;
        RECT 40.105 2704.755 40.395 2704.800 ;
        RECT 41.010 2704.740 41.330 2704.800 ;
        RECT 41.010 2608.380 41.330 2608.440 ;
        RECT 41.930 2608.380 42.250 2608.440 ;
        RECT 41.010 2608.240 42.250 2608.380 ;
        RECT 41.010 2608.180 41.330 2608.240 ;
        RECT 41.930 2608.180 42.250 2608.240 ;
        RECT 41.010 2511.820 41.330 2511.880 ;
        RECT 41.930 2511.820 42.250 2511.880 ;
        RECT 41.010 2511.680 42.250 2511.820 ;
        RECT 41.010 2511.620 41.330 2511.680 ;
        RECT 41.930 2511.620 42.250 2511.680 ;
        RECT 39.630 2463.200 39.950 2463.260 ;
        RECT 40.550 2463.200 40.870 2463.260 ;
        RECT 39.630 2463.060 40.870 2463.200 ;
        RECT 39.630 2463.000 39.950 2463.060 ;
        RECT 40.550 2463.000 40.870 2463.060 ;
        RECT 40.090 2366.640 40.410 2366.700 ;
        RECT 40.550 2366.640 40.870 2366.700 ;
        RECT 40.090 2366.500 40.870 2366.640 ;
        RECT 40.090 2366.440 40.410 2366.500 ;
        RECT 40.550 2366.440 40.870 2366.500 ;
        RECT 40.090 2235.540 40.410 2235.800 ;
        RECT 40.180 2235.400 40.320 2235.540 ;
        RECT 40.550 2235.400 40.870 2235.460 ;
        RECT 40.180 2235.260 40.870 2235.400 ;
        RECT 40.550 2235.200 40.870 2235.260 ;
        RECT 39.170 2221.800 39.490 2221.860 ;
        RECT 40.550 2221.800 40.870 2221.860 ;
        RECT 39.170 2221.660 40.870 2221.800 ;
        RECT 39.170 2221.600 39.490 2221.660 ;
        RECT 40.550 2221.600 40.870 2221.660 ;
        RECT 40.090 2139.320 40.410 2139.580 ;
        RECT 40.180 2138.900 40.320 2139.320 ;
        RECT 40.090 2138.640 40.410 2138.900 ;
        RECT 40.090 2090.900 40.410 2090.960 ;
        RECT 41.010 2090.900 41.330 2090.960 ;
        RECT 40.090 2090.760 41.330 2090.900 ;
        RECT 40.090 2090.700 40.410 2090.760 ;
        RECT 41.010 2090.700 41.330 2090.760 ;
        RECT 40.090 1994.680 40.410 1994.740 ;
        RECT 39.895 1994.540 40.410 1994.680 ;
        RECT 40.090 1994.480 40.410 1994.540 ;
        RECT 40.090 1952.860 40.410 1952.920 ;
        RECT 39.895 1952.720 40.410 1952.860 ;
        RECT 40.090 1952.660 40.410 1952.720 ;
        RECT 39.170 1904.580 39.490 1904.640 ;
        RECT 40.090 1904.580 40.410 1904.640 ;
        RECT 39.170 1904.440 40.410 1904.580 ;
        RECT 39.170 1904.380 39.490 1904.440 ;
        RECT 40.090 1904.380 40.410 1904.440 ;
        RECT 40.090 1849.500 40.410 1849.560 ;
        RECT 39.720 1849.360 40.410 1849.500 ;
        RECT 39.720 1849.220 39.860 1849.360 ;
        RECT 40.090 1849.300 40.410 1849.360 ;
        RECT 39.630 1848.960 39.950 1849.220 ;
        RECT 39.630 1800.880 39.950 1800.940 ;
        RECT 40.550 1800.880 40.870 1800.940 ;
        RECT 39.630 1800.740 40.870 1800.880 ;
        RECT 39.630 1800.680 39.950 1800.740 ;
        RECT 40.550 1800.680 40.870 1800.740 ;
        RECT 40.105 1786.940 40.395 1786.985 ;
        RECT 40.550 1786.940 40.870 1787.000 ;
        RECT 40.105 1786.800 40.870 1786.940 ;
        RECT 40.105 1786.755 40.395 1786.800 ;
        RECT 40.550 1786.740 40.870 1786.800 ;
        RECT 40.090 1739.000 40.410 1739.060 ;
        RECT 39.895 1738.860 40.410 1739.000 ;
        RECT 40.090 1738.800 40.410 1738.860 ;
        RECT 40.090 1705.000 40.410 1705.060 ;
        RECT 39.895 1704.860 40.410 1705.000 ;
        RECT 40.090 1704.800 40.410 1704.860 ;
        RECT 40.090 1684.260 40.410 1684.320 ;
        RECT 39.895 1684.120 40.410 1684.260 ;
        RECT 40.090 1684.060 40.410 1684.120 ;
        RECT 39.645 1683.240 39.935 1683.285 ;
        RECT 40.090 1683.240 40.410 1683.300 ;
        RECT 39.645 1683.100 40.410 1683.240 ;
        RECT 39.645 1683.055 39.935 1683.100 ;
        RECT 40.090 1683.040 40.410 1683.100 ;
        RECT 39.630 1635.640 39.950 1635.700 ;
        RECT 39.435 1635.500 39.950 1635.640 ;
        RECT 39.630 1635.440 39.950 1635.500 ;
        RECT 39.630 1607.420 39.950 1607.480 ;
        RECT 41.010 1607.420 41.330 1607.480 ;
        RECT 39.630 1607.280 41.330 1607.420 ;
        RECT 39.630 1607.220 39.950 1607.280 ;
        RECT 41.010 1607.220 41.330 1607.280 ;
        RECT 39.630 1546.220 39.950 1546.280 ;
        RECT 41.010 1546.220 41.330 1546.280 ;
        RECT 39.630 1546.080 41.330 1546.220 ;
        RECT 39.630 1546.020 39.950 1546.080 ;
        RECT 41.010 1546.020 41.330 1546.080 ;
        RECT 40.090 1511.340 40.410 1511.600 ;
        RECT 40.180 1510.520 40.320 1511.340 ;
        RECT 40.550 1510.520 40.870 1510.580 ;
        RECT 40.180 1510.380 40.870 1510.520 ;
        RECT 40.550 1510.320 40.870 1510.380 ;
        RECT 40.565 1448.980 40.855 1449.025 ;
        RECT 41.010 1448.980 41.330 1449.040 ;
        RECT 40.565 1448.840 41.330 1448.980 ;
        RECT 40.565 1448.795 40.855 1448.840 ;
        RECT 41.010 1448.780 41.330 1448.840 ;
        RECT 40.550 1401.040 40.870 1401.100 ;
        RECT 40.355 1400.900 40.870 1401.040 ;
        RECT 40.550 1400.840 40.870 1400.900 ;
        RECT 40.550 1366.500 40.870 1366.760 ;
        RECT 40.640 1365.740 40.780 1366.500 ;
        RECT 40.550 1365.480 40.870 1365.740 ;
        RECT 39.630 1159.300 39.950 1159.360 ;
        RECT 40.090 1159.300 40.410 1159.360 ;
        RECT 39.630 1159.160 40.410 1159.300 ;
        RECT 39.630 1159.100 39.950 1159.160 ;
        RECT 40.090 1159.100 40.410 1159.160 ;
        RECT 40.090 1110.680 40.410 1110.740 ;
        RECT 39.895 1110.540 40.410 1110.680 ;
        RECT 40.090 1110.480 40.410 1110.540 ;
        RECT 40.105 1076.000 40.395 1076.045 ;
        RECT 40.550 1076.000 40.870 1076.060 ;
        RECT 40.105 1075.860 40.870 1076.000 ;
        RECT 40.105 1075.815 40.395 1075.860 ;
        RECT 40.550 1075.800 40.870 1075.860 ;
        RECT 40.550 1028.740 40.870 1028.800 ;
        RECT 39.720 1028.600 40.870 1028.740 ;
        RECT 39.720 1028.120 39.860 1028.600 ;
        RECT 40.550 1028.540 40.870 1028.600 ;
        RECT 39.630 1027.860 39.950 1028.120 ;
        RECT 39.630 1007.320 39.950 1007.380 ;
        RECT 39.435 1007.180 39.950 1007.320 ;
        RECT 39.630 1007.120 39.950 1007.180 ;
        RECT 39.630 965.840 39.950 965.900 ;
        RECT 39.435 965.700 39.950 965.840 ;
        RECT 39.630 965.640 39.950 965.700 ;
        RECT 40.090 931.840 40.410 931.900 ;
        RECT 40.090 931.700 40.780 931.840 ;
        RECT 40.090 931.640 40.410 931.700 ;
        RECT 40.640 931.220 40.780 931.700 ;
        RECT 40.550 930.960 40.870 931.220 ;
        RECT 40.550 883.700 40.870 883.960 ;
        RECT 40.090 882.880 40.410 882.940 ;
        RECT 40.640 882.880 40.780 883.700 ;
        RECT 40.090 882.740 40.780 882.880 ;
        RECT 40.090 882.680 40.410 882.740 ;
        RECT 40.090 821.000 40.410 821.060 ;
        RECT 40.550 821.000 40.870 821.060 ;
        RECT 40.090 820.860 40.870 821.000 ;
        RECT 40.090 820.800 40.410 820.860 ;
        RECT 40.550 820.800 40.870 820.860 ;
        RECT 40.090 724.440 40.410 724.500 ;
        RECT 40.550 724.440 40.870 724.500 ;
        RECT 40.090 724.300 40.870 724.440 ;
        RECT 40.090 724.240 40.410 724.300 ;
        RECT 40.550 724.240 40.870 724.300 ;
        RECT 39.645 627.880 39.935 627.925 ;
        RECT 40.090 627.880 40.410 627.940 ;
        RECT 39.645 627.740 40.410 627.880 ;
        RECT 39.645 627.695 39.935 627.740 ;
        RECT 40.090 627.680 40.410 627.740 ;
        RECT 39.630 579.940 39.950 580.000 ;
        RECT 39.435 579.800 39.950 579.940 ;
        RECT 39.630 579.740 39.950 579.800 ;
        RECT 40.090 531.320 40.410 531.380 ;
        RECT 39.895 531.180 40.410 531.320 ;
        RECT 40.090 531.120 40.410 531.180 ;
        RECT 40.090 496.640 40.410 496.700 ;
        RECT 39.895 496.500 40.410 496.640 ;
        RECT 40.090 496.440 40.410 496.500 ;
        RECT 40.550 455.160 40.870 455.220 ;
        RECT 296.770 455.160 297.090 455.220 ;
        RECT 40.550 455.020 297.090 455.160 ;
        RECT 40.550 454.960 40.870 455.020 ;
        RECT 296.770 454.960 297.090 455.020 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3270.500 40.380 3270.760 ;
        RECT 41.040 3270.500 41.300 3270.760 ;
        RECT 40.120 3173.940 40.380 3174.200 ;
        RECT 41.040 3173.940 41.300 3174.200 ;
        RECT 40.120 3077.380 40.380 3077.640 ;
        RECT 41.040 3077.380 41.300 3077.640 ;
        RECT 40.120 2980.820 40.380 2981.080 ;
        RECT 41.040 2980.820 41.300 2981.080 ;
        RECT 40.120 2946.140 40.380 2946.400 ;
        RECT 40.120 2898.540 40.380 2898.800 ;
        RECT 39.660 2897.860 39.920 2898.120 ;
        RECT 40.580 2897.860 40.840 2898.120 ;
        RECT 39.660 2814.560 39.920 2814.820 ;
        RECT 40.580 2814.560 40.840 2814.820 ;
        RECT 40.120 2752.680 40.380 2752.940 ;
        RECT 41.040 2704.740 41.300 2705.000 ;
        RECT 41.040 2608.180 41.300 2608.440 ;
        RECT 41.960 2608.180 42.220 2608.440 ;
        RECT 41.040 2511.620 41.300 2511.880 ;
        RECT 41.960 2511.620 42.220 2511.880 ;
        RECT 39.660 2463.000 39.920 2463.260 ;
        RECT 40.580 2463.000 40.840 2463.260 ;
        RECT 40.120 2366.440 40.380 2366.700 ;
        RECT 40.580 2366.440 40.840 2366.700 ;
        RECT 40.120 2235.540 40.380 2235.800 ;
        RECT 40.580 2235.200 40.840 2235.460 ;
        RECT 39.200 2221.600 39.460 2221.860 ;
        RECT 40.580 2221.600 40.840 2221.860 ;
        RECT 40.120 2139.320 40.380 2139.580 ;
        RECT 40.120 2138.640 40.380 2138.900 ;
        RECT 40.120 2090.700 40.380 2090.960 ;
        RECT 41.040 2090.700 41.300 2090.960 ;
        RECT 40.120 1994.480 40.380 1994.740 ;
        RECT 40.120 1952.660 40.380 1952.920 ;
        RECT 39.200 1904.380 39.460 1904.640 ;
        RECT 40.120 1904.380 40.380 1904.640 ;
        RECT 40.120 1849.300 40.380 1849.560 ;
        RECT 39.660 1848.960 39.920 1849.220 ;
        RECT 39.660 1800.680 39.920 1800.940 ;
        RECT 40.580 1800.680 40.840 1800.940 ;
        RECT 40.580 1786.740 40.840 1787.000 ;
        RECT 40.120 1738.800 40.380 1739.060 ;
        RECT 40.120 1704.800 40.380 1705.060 ;
        RECT 40.120 1684.060 40.380 1684.320 ;
        RECT 40.120 1683.040 40.380 1683.300 ;
        RECT 39.660 1635.440 39.920 1635.700 ;
        RECT 39.660 1607.220 39.920 1607.480 ;
        RECT 41.040 1607.220 41.300 1607.480 ;
        RECT 39.660 1546.020 39.920 1546.280 ;
        RECT 41.040 1546.020 41.300 1546.280 ;
        RECT 40.120 1511.340 40.380 1511.600 ;
        RECT 40.580 1510.320 40.840 1510.580 ;
        RECT 41.040 1448.780 41.300 1449.040 ;
        RECT 40.580 1400.840 40.840 1401.100 ;
        RECT 40.580 1366.500 40.840 1366.760 ;
        RECT 40.580 1365.480 40.840 1365.740 ;
        RECT 39.660 1159.100 39.920 1159.360 ;
        RECT 40.120 1159.100 40.380 1159.360 ;
        RECT 40.120 1110.480 40.380 1110.740 ;
        RECT 40.580 1075.800 40.840 1076.060 ;
        RECT 40.580 1028.540 40.840 1028.800 ;
        RECT 39.660 1027.860 39.920 1028.120 ;
        RECT 39.660 1007.120 39.920 1007.380 ;
        RECT 39.660 965.640 39.920 965.900 ;
        RECT 40.120 931.640 40.380 931.900 ;
        RECT 40.580 930.960 40.840 931.220 ;
        RECT 40.580 883.700 40.840 883.960 ;
        RECT 40.120 882.680 40.380 882.940 ;
        RECT 40.120 820.800 40.380 821.060 ;
        RECT 40.580 820.800 40.840 821.060 ;
        RECT 40.120 724.240 40.380 724.500 ;
        RECT 40.580 724.240 40.840 724.500 ;
        RECT 40.120 627.680 40.380 627.940 ;
        RECT 39.660 579.740 39.920 580.000 ;
        RECT 40.120 531.120 40.380 531.380 ;
        RECT 40.120 496.440 40.380 496.700 ;
        RECT 40.580 454.960 40.840 455.220 ;
        RECT 296.800 454.960 297.060 455.220 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3270.790 40.320 3318.670 ;
        RECT 40.120 3270.470 40.380 3270.790 ;
        RECT 41.040 3270.470 41.300 3270.790 ;
        RECT 41.100 3222.250 41.240 3270.470 ;
        RECT 40.180 3222.110 41.240 3222.250 ;
        RECT 40.180 3174.230 40.320 3222.110 ;
        RECT 40.120 3173.910 40.380 3174.230 ;
        RECT 41.040 3173.910 41.300 3174.230 ;
        RECT 41.100 3125.690 41.240 3173.910 ;
        RECT 40.180 3125.550 41.240 3125.690 ;
        RECT 40.180 3077.670 40.320 3125.550 ;
        RECT 40.120 3077.350 40.380 3077.670 ;
        RECT 41.040 3077.350 41.300 3077.670 ;
        RECT 41.100 3029.130 41.240 3077.350 ;
        RECT 40.180 3028.990 41.240 3029.130 ;
        RECT 40.180 2981.110 40.320 3028.990 ;
        RECT 40.120 2980.790 40.380 2981.110 ;
        RECT 41.040 2980.850 41.300 2981.110 ;
        RECT 40.640 2980.790 41.300 2980.850 ;
        RECT 40.640 2980.710 41.240 2980.790 ;
        RECT 40.640 2959.770 40.780 2980.710 ;
        RECT 40.180 2959.630 40.780 2959.770 ;
        RECT 40.180 2946.430 40.320 2959.630 ;
        RECT 40.120 2946.110 40.380 2946.430 ;
        RECT 40.120 2898.570 40.380 2898.830 ;
        RECT 39.720 2898.510 40.380 2898.570 ;
        RECT 39.720 2898.430 40.320 2898.510 ;
        RECT 39.720 2898.150 39.860 2898.430 ;
        RECT 39.660 2897.830 39.920 2898.150 ;
        RECT 40.580 2897.830 40.840 2898.150 ;
        RECT 40.640 2814.850 40.780 2897.830 ;
        RECT 39.660 2814.530 39.920 2814.850 ;
        RECT 40.580 2814.530 40.840 2814.850 ;
        RECT 39.720 2766.650 39.860 2814.530 ;
        RECT 39.720 2766.510 40.320 2766.650 ;
        RECT 40.180 2752.970 40.320 2766.510 ;
        RECT 40.120 2752.650 40.380 2752.970 ;
        RECT 41.040 2704.710 41.300 2705.030 ;
        RECT 41.100 2670.090 41.240 2704.710 ;
        RECT 40.640 2669.950 41.240 2670.090 ;
        RECT 40.640 2656.605 40.780 2669.950 ;
        RECT 40.570 2656.235 40.850 2656.605 ;
        RECT 41.950 2656.235 42.230 2656.605 ;
        RECT 42.020 2608.470 42.160 2656.235 ;
        RECT 41.040 2608.150 41.300 2608.470 ;
        RECT 41.960 2608.150 42.220 2608.470 ;
        RECT 41.100 2573.530 41.240 2608.150 ;
        RECT 40.640 2573.390 41.240 2573.530 ;
        RECT 40.640 2560.045 40.780 2573.390 ;
        RECT 40.570 2559.675 40.850 2560.045 ;
        RECT 41.950 2559.675 42.230 2560.045 ;
        RECT 42.020 2511.910 42.160 2559.675 ;
        RECT 41.040 2511.590 41.300 2511.910 ;
        RECT 41.960 2511.590 42.220 2511.910 ;
        RECT 41.100 2476.970 41.240 2511.590 ;
        RECT 40.640 2476.830 41.240 2476.970 ;
        RECT 40.640 2463.290 40.780 2476.830 ;
        RECT 39.660 2462.970 39.920 2463.290 ;
        RECT 40.580 2462.970 40.840 2463.290 ;
        RECT 39.720 2415.205 39.860 2462.970 ;
        RECT 39.650 2414.835 39.930 2415.205 ;
        RECT 41.030 2414.835 41.310 2415.205 ;
        RECT 41.100 2380.410 41.240 2414.835 ;
        RECT 40.180 2380.270 41.240 2380.410 ;
        RECT 40.180 2366.730 40.320 2380.270 ;
        RECT 40.120 2366.410 40.380 2366.730 ;
        RECT 40.580 2366.410 40.840 2366.730 ;
        RECT 40.640 2318.530 40.780 2366.410 ;
        RECT 40.640 2318.390 41.240 2318.530 ;
        RECT 41.100 2283.850 41.240 2318.390 ;
        RECT 40.180 2283.710 41.240 2283.850 ;
        RECT 40.180 2235.830 40.320 2283.710 ;
        RECT 40.120 2235.510 40.380 2235.830 ;
        RECT 40.580 2235.170 40.840 2235.490 ;
        RECT 40.640 2221.890 40.780 2235.170 ;
        RECT 39.200 2221.570 39.460 2221.890 ;
        RECT 40.580 2221.570 40.840 2221.890 ;
        RECT 39.260 2173.805 39.400 2221.570 ;
        RECT 39.190 2173.435 39.470 2173.805 ;
        RECT 40.110 2173.435 40.390 2173.805 ;
        RECT 40.180 2139.610 40.320 2173.435 ;
        RECT 40.120 2139.290 40.380 2139.610 ;
        RECT 40.120 2138.610 40.380 2138.930 ;
        RECT 40.180 2090.990 40.320 2138.610 ;
        RECT 40.120 2090.670 40.380 2090.990 ;
        RECT 41.040 2090.670 41.300 2090.990 ;
        RECT 41.100 2042.450 41.240 2090.670 ;
        RECT 40.180 2042.310 41.240 2042.450 ;
        RECT 40.180 1994.770 40.320 2042.310 ;
        RECT 40.120 1994.450 40.380 1994.770 ;
        RECT 40.180 1952.950 40.320 1953.105 ;
        RECT 40.120 1952.690 40.380 1952.950 ;
        RECT 39.260 1952.630 40.380 1952.690 ;
        RECT 39.260 1952.550 40.320 1952.630 ;
        RECT 39.260 1904.670 39.400 1952.550 ;
        RECT 39.200 1904.350 39.460 1904.670 ;
        RECT 40.120 1904.350 40.380 1904.670 ;
        RECT 40.180 1849.590 40.320 1904.350 ;
        RECT 40.120 1849.270 40.380 1849.590 ;
        RECT 39.660 1848.930 39.920 1849.250 ;
        RECT 39.720 1800.970 39.860 1848.930 ;
        RECT 39.660 1800.650 39.920 1800.970 ;
        RECT 40.580 1800.650 40.840 1800.970 ;
        RECT 40.640 1787.030 40.780 1800.650 ;
        RECT 40.580 1786.710 40.840 1787.030 ;
        RECT 40.120 1738.770 40.380 1739.090 ;
        RECT 40.180 1705.090 40.320 1738.770 ;
        RECT 40.120 1704.770 40.380 1705.090 ;
        RECT 40.120 1684.030 40.380 1684.350 ;
        RECT 40.180 1683.330 40.320 1684.030 ;
        RECT 40.120 1683.010 40.380 1683.330 ;
        RECT 39.660 1635.410 39.920 1635.730 ;
        RECT 39.720 1607.510 39.860 1635.410 ;
        RECT 39.660 1607.190 39.920 1607.510 ;
        RECT 41.040 1607.190 41.300 1607.510 ;
        RECT 41.100 1546.310 41.240 1607.190 ;
        RECT 39.660 1546.050 39.920 1546.310 ;
        RECT 39.660 1545.990 40.320 1546.050 ;
        RECT 41.040 1545.990 41.300 1546.310 ;
        RECT 39.720 1545.910 40.320 1545.990 ;
        RECT 40.180 1511.630 40.320 1545.910 ;
        RECT 40.120 1511.310 40.380 1511.630 ;
        RECT 40.580 1510.290 40.840 1510.610 ;
        RECT 40.640 1463.090 40.780 1510.290 ;
        RECT 40.640 1462.950 41.240 1463.090 ;
        RECT 41.100 1449.070 41.240 1462.950 ;
        RECT 41.040 1448.750 41.300 1449.070 ;
        RECT 40.580 1400.810 40.840 1401.130 ;
        RECT 40.640 1366.790 40.780 1400.810 ;
        RECT 40.580 1366.470 40.840 1366.790 ;
        RECT 40.580 1365.450 40.840 1365.770 ;
        RECT 40.640 1221.010 40.780 1365.450 ;
        RECT 40.180 1220.870 40.780 1221.010 ;
        RECT 40.180 1159.390 40.320 1220.870 ;
        RECT 39.660 1159.070 39.920 1159.390 ;
        RECT 40.120 1159.070 40.380 1159.390 ;
        RECT 39.720 1124.450 39.860 1159.070 ;
        RECT 39.720 1124.310 40.320 1124.450 ;
        RECT 40.180 1110.770 40.320 1124.310 ;
        RECT 40.120 1110.450 40.380 1110.770 ;
        RECT 40.580 1075.770 40.840 1076.090 ;
        RECT 40.640 1028.830 40.780 1075.770 ;
        RECT 40.580 1028.510 40.840 1028.830 ;
        RECT 39.660 1027.830 39.920 1028.150 ;
        RECT 39.720 1007.410 39.860 1027.830 ;
        RECT 39.660 1007.090 39.920 1007.410 ;
        RECT 39.660 965.610 39.920 965.930 ;
        RECT 39.720 959.210 39.860 965.610 ;
        RECT 39.720 959.070 40.320 959.210 ;
        RECT 40.180 931.930 40.320 959.070 ;
        RECT 40.120 931.610 40.380 931.930 ;
        RECT 40.580 930.930 40.840 931.250 ;
        RECT 40.640 883.990 40.780 930.930 ;
        RECT 40.580 883.670 40.840 883.990 ;
        RECT 40.120 882.650 40.380 882.970 ;
        RECT 40.180 821.090 40.320 882.650 ;
        RECT 40.120 820.770 40.380 821.090 ;
        RECT 40.580 820.770 40.840 821.090 ;
        RECT 40.640 772.890 40.780 820.770 ;
        RECT 40.640 772.750 41.240 772.890 ;
        RECT 41.100 738.210 41.240 772.750 ;
        RECT 40.180 738.070 41.240 738.210 ;
        RECT 40.180 724.530 40.320 738.070 ;
        RECT 40.120 724.210 40.380 724.530 ;
        RECT 40.580 724.210 40.840 724.530 ;
        RECT 40.640 676.330 40.780 724.210 ;
        RECT 40.640 676.190 41.240 676.330 ;
        RECT 41.100 641.650 41.240 676.190 ;
        RECT 40.180 641.510 41.240 641.650 ;
        RECT 40.180 627.970 40.320 641.510 ;
        RECT 40.120 627.650 40.380 627.970 ;
        RECT 39.660 579.710 39.920 580.030 ;
        RECT 39.720 545.090 39.860 579.710 ;
        RECT 39.720 544.950 40.320 545.090 ;
        RECT 40.180 531.410 40.320 544.950 ;
        RECT 40.120 531.090 40.380 531.410 ;
        RECT 40.120 496.410 40.380 496.730 ;
        RECT 40.180 483.210 40.320 496.410 ;
        RECT 40.180 483.070 40.780 483.210 ;
        RECT 40.640 455.250 40.780 483.070 ;
        RECT 40.580 454.930 40.840 455.250 ;
        RECT 296.800 454.930 297.060 455.250 ;
        RECT 296.860 454.765 297.000 454.930 ;
        RECT 296.790 454.395 297.070 454.765 ;
      LAYER via2 ;
        RECT 40.570 2656.280 40.850 2656.560 ;
        RECT 41.950 2656.280 42.230 2656.560 ;
        RECT 40.570 2559.720 40.850 2560.000 ;
        RECT 41.950 2559.720 42.230 2560.000 ;
        RECT 39.650 2414.880 39.930 2415.160 ;
        RECT 41.030 2414.880 41.310 2415.160 ;
        RECT 39.190 2173.480 39.470 2173.760 ;
        RECT 40.110 2173.480 40.390 2173.760 ;
        RECT 296.790 454.440 297.070 454.720 ;
      LAYER met3 ;
        RECT 40.545 2656.570 40.875 2656.585 ;
        RECT 41.925 2656.570 42.255 2656.585 ;
        RECT 40.545 2656.270 42.255 2656.570 ;
        RECT 40.545 2656.255 40.875 2656.270 ;
        RECT 41.925 2656.255 42.255 2656.270 ;
        RECT 40.545 2560.010 40.875 2560.025 ;
        RECT 41.925 2560.010 42.255 2560.025 ;
        RECT 40.545 2559.710 42.255 2560.010 ;
        RECT 40.545 2559.695 40.875 2559.710 ;
        RECT 41.925 2559.695 42.255 2559.710 ;
        RECT 39.625 2415.170 39.955 2415.185 ;
        RECT 41.005 2415.170 41.335 2415.185 ;
        RECT 39.625 2414.870 41.335 2415.170 ;
        RECT 39.625 2414.855 39.955 2414.870 ;
        RECT 41.005 2414.855 41.335 2414.870 ;
        RECT 39.165 2173.770 39.495 2173.785 ;
        RECT 40.085 2173.770 40.415 2173.785 ;
        RECT 39.165 2173.470 40.415 2173.770 ;
        RECT 39.165 2173.455 39.495 2173.470 ;
        RECT 40.085 2173.455 40.415 2173.470 ;
        RECT 296.765 454.730 297.095 454.745 ;
        RECT 296.765 454.640 310.500 454.730 ;
        RECT 296.765 454.430 314.000 454.640 ;
        RECT 296.765 454.415 297.095 454.430 ;
        RECT 310.000 454.040 314.000 454.430 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 3267.555 16.930 3267.925 ;
        RECT 16.720 3264.525 16.860 3267.555 ;
        RECT 16.650 3264.155 16.930 3264.525 ;
        RECT 792.170 216.000 792.450 220.000 ;
        RECT 792.280 212.685 792.420 216.000 ;
        RECT 792.210 212.315 792.490 212.685 ;
      LAYER via2 ;
        RECT 16.650 3267.600 16.930 3267.880 ;
        RECT 16.650 3264.200 16.930 3264.480 ;
        RECT 792.210 212.360 792.490 212.640 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 16.625 3267.890 16.955 3267.905 ;
        RECT -4.800 3267.590 16.955 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 16.625 3267.575 16.955 3267.590 ;
        RECT 16.625 3264.490 16.955 3264.505 ;
        RECT 285.470 3264.490 285.850 3264.500 ;
        RECT 16.625 3264.190 285.850 3264.490 ;
        RECT 16.625 3264.175 16.955 3264.190 ;
        RECT 285.470 3264.180 285.850 3264.190 ;
        RECT 285.470 212.650 285.850 212.660 ;
        RECT 792.185 212.650 792.515 212.665 ;
        RECT 285.470 212.350 792.515 212.650 ;
        RECT 285.470 212.340 285.850 212.350 ;
        RECT 792.185 212.335 792.515 212.350 ;
      LAYER via3 ;
        RECT 285.500 3264.180 285.820 3264.500 ;
        RECT 285.500 212.340 285.820 212.660 ;
      LAYER met4 ;
        RECT 285.495 3264.175 285.825 3264.505 ;
        RECT 285.510 212.665 285.810 3264.175 ;
        RECT 285.495 212.335 285.825 212.665 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 2974.220 16.490 2974.280 ;
        RECT 952.270 2974.220 952.590 2974.280 ;
        RECT 16.170 2974.080 952.590 2974.220 ;
        RECT 16.170 2974.020 16.490 2974.080 ;
        RECT 952.270 2974.020 952.590 2974.080 ;
      LAYER via ;
        RECT 16.200 2974.020 16.460 2974.280 ;
        RECT 952.300 2974.020 952.560 2974.280 ;
      LAYER met2 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 16.260 2974.310 16.400 2979.915 ;
        RECT 16.200 2973.990 16.460 2974.310 ;
        RECT 952.300 2973.990 952.560 2974.310 ;
        RECT 952.360 1325.730 952.500 2973.990 ;
        RECT 952.360 1325.590 954.800 1325.730 ;
        RECT 954.660 1324.370 954.800 1325.590 ;
        RECT 957.770 1324.370 958.050 1325.025 ;
        RECT 954.660 1324.230 958.050 1324.370 ;
        RECT 957.770 1321.025 958.050 1324.230 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.800 2979.950 16.495 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 19.850 2692.360 20.170 2692.420 ;
        RECT 51.590 2692.360 51.910 2692.420 ;
        RECT 19.850 2692.220 51.910 2692.360 ;
        RECT 19.850 2692.160 20.170 2692.220 ;
        RECT 51.590 2692.160 51.910 2692.220 ;
        RECT 51.590 393.280 51.910 393.340 ;
        RECT 296.770 393.280 297.090 393.340 ;
        RECT 51.590 393.140 297.090 393.280 ;
        RECT 51.590 393.080 51.910 393.140 ;
        RECT 296.770 393.080 297.090 393.140 ;
      LAYER via ;
        RECT 19.880 2692.160 20.140 2692.420 ;
        RECT 51.620 2692.160 51.880 2692.420 ;
        RECT 51.620 393.080 51.880 393.340 ;
        RECT 296.800 393.080 297.060 393.340 ;
      LAYER met2 ;
        RECT 19.870 2692.955 20.150 2693.325 ;
        RECT 19.940 2692.450 20.080 2692.955 ;
        RECT 19.880 2692.130 20.140 2692.450 ;
        RECT 51.620 2692.130 51.880 2692.450 ;
        RECT 51.680 393.370 51.820 2692.130 ;
        RECT 51.620 393.050 51.880 393.370 ;
        RECT 296.800 393.050 297.060 393.370 ;
        RECT 296.860 388.125 297.000 393.050 ;
        RECT 296.790 387.755 297.070 388.125 ;
      LAYER via2 ;
        RECT 19.870 2693.000 20.150 2693.280 ;
        RECT 296.790 387.800 297.070 388.080 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 19.845 2693.290 20.175 2693.305 ;
        RECT -4.800 2692.990 20.175 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 19.845 2692.975 20.175 2692.990 ;
        RECT 296.765 388.090 297.095 388.105 ;
        RECT 296.765 388.000 310.500 388.090 ;
        RECT 296.765 387.790 314.000 388.000 ;
        RECT 296.765 387.775 297.095 387.790 ;
        RECT 310.000 387.400 314.000 387.790 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2403.020 16.950 2403.080 ;
        RECT 58.490 2403.020 58.810 2403.080 ;
        RECT 16.630 2402.880 58.810 2403.020 ;
        RECT 16.630 2402.820 16.950 2402.880 ;
        RECT 58.490 2402.820 58.810 2402.880 ;
        RECT 58.490 205.600 58.810 205.660 ;
        RECT 446.270 205.600 446.590 205.660 ;
        RECT 58.490 205.460 446.590 205.600 ;
        RECT 58.490 205.400 58.810 205.460 ;
        RECT 446.270 205.400 446.590 205.460 ;
      LAYER via ;
        RECT 16.660 2402.820 16.920 2403.080 ;
        RECT 58.520 2402.820 58.780 2403.080 ;
        RECT 58.520 205.400 58.780 205.660 ;
        RECT 446.300 205.400 446.560 205.660 ;
      LAYER met2 ;
        RECT 16.650 2405.315 16.930 2405.685 ;
        RECT 16.720 2403.110 16.860 2405.315 ;
        RECT 16.660 2402.790 16.920 2403.110 ;
        RECT 58.520 2402.790 58.780 2403.110 ;
        RECT 58.580 205.690 58.720 2402.790 ;
        RECT 446.250 216.000 446.530 220.000 ;
        RECT 446.360 205.690 446.500 216.000 ;
        RECT 58.520 205.370 58.780 205.690 ;
        RECT 446.300 205.370 446.560 205.690 ;
      LAYER via2 ;
        RECT 16.650 2405.360 16.930 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 16.625 2405.650 16.955 2405.665 ;
        RECT -4.800 2405.350 16.955 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 16.625 2405.335 16.955 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 2118.440 20.630 2118.500 ;
        RECT 65.390 2118.440 65.710 2118.500 ;
        RECT 20.310 2118.300 65.710 2118.440 ;
        RECT 20.310 2118.240 20.630 2118.300 ;
        RECT 65.390 2118.240 65.710 2118.300 ;
        RECT 65.390 827.800 65.710 827.860 ;
        RECT 296.770 827.800 297.090 827.860 ;
        RECT 65.390 827.660 297.090 827.800 ;
        RECT 65.390 827.600 65.710 827.660 ;
        RECT 296.770 827.600 297.090 827.660 ;
      LAYER via ;
        RECT 20.340 2118.240 20.600 2118.500 ;
        RECT 65.420 2118.240 65.680 2118.500 ;
        RECT 65.420 827.600 65.680 827.860 ;
        RECT 296.800 827.600 297.060 827.860 ;
      LAYER met2 ;
        RECT 20.330 2118.355 20.610 2118.725 ;
        RECT 20.340 2118.210 20.600 2118.355 ;
        RECT 65.420 2118.210 65.680 2118.530 ;
        RECT 65.480 827.890 65.620 2118.210 ;
        RECT 65.420 827.570 65.680 827.890 ;
        RECT 296.800 827.570 297.060 827.890 ;
        RECT 296.860 827.405 297.000 827.570 ;
        RECT 296.790 827.035 297.070 827.405 ;
      LAYER via2 ;
        RECT 20.330 2118.400 20.610 2118.680 ;
        RECT 296.790 827.080 297.070 827.360 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 20.305 2118.690 20.635 2118.705 ;
        RECT -4.800 2118.390 20.635 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 20.305 2118.375 20.635 2118.390 ;
        RECT 296.765 827.370 297.095 827.385 ;
        RECT 296.765 827.280 310.500 827.370 ;
        RECT 296.765 827.070 314.000 827.280 ;
        RECT 296.765 827.055 297.095 827.070 ;
        RECT 310.000 826.680 314.000 827.070 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 1828.760 20.630 1828.820 ;
        RECT 917.770 1828.760 918.090 1828.820 ;
        RECT 20.310 1828.620 918.090 1828.760 ;
        RECT 20.310 1828.560 20.630 1828.620 ;
        RECT 917.770 1828.560 918.090 1828.620 ;
      LAYER via ;
        RECT 20.340 1828.560 20.600 1828.820 ;
        RECT 917.800 1828.560 918.060 1828.820 ;
      LAYER met2 ;
        RECT 20.330 1830.715 20.610 1831.085 ;
        RECT 20.400 1828.850 20.540 1830.715 ;
        RECT 20.340 1828.530 20.600 1828.850 ;
        RECT 917.800 1828.530 918.060 1828.850 ;
        RECT 917.860 1325.050 918.000 1828.530 ;
        RECT 917.860 1325.025 918.390 1325.050 ;
        RECT 917.860 1324.910 918.490 1325.025 ;
        RECT 918.210 1321.025 918.490 1324.910 ;
      LAYER via2 ;
        RECT 20.330 1830.760 20.610 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 20.305 1831.050 20.635 1831.065 ;
        RECT -4.800 1830.750 20.635 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 20.305 1830.735 20.635 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1542.450 669.700 1542.770 669.760 ;
        RECT 2900.830 669.700 2901.150 669.760 ;
        RECT 1542.450 669.560 2901.150 669.700 ;
        RECT 1542.450 669.500 1542.770 669.560 ;
        RECT 2900.830 669.500 2901.150 669.560 ;
        RECT 1419.170 448.360 1419.490 448.420 ;
        RECT 1542.450 448.360 1542.770 448.420 ;
        RECT 1419.170 448.220 1542.770 448.360 ;
        RECT 1419.170 448.160 1419.490 448.220 ;
        RECT 1542.450 448.160 1542.770 448.220 ;
      LAYER via ;
        RECT 1542.480 669.500 1542.740 669.760 ;
        RECT 2900.860 669.500 2901.120 669.760 ;
        RECT 1419.200 448.160 1419.460 448.420 ;
        RECT 1542.480 448.160 1542.740 448.420 ;
      LAYER met2 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
        RECT 2900.920 669.790 2901.060 674.035 ;
        RECT 1542.480 669.470 1542.740 669.790 ;
        RECT 2900.860 669.470 2901.120 669.790 ;
        RECT 1542.540 448.450 1542.680 669.470 ;
        RECT 1419.200 448.130 1419.460 448.450 ;
        RECT 1542.480 448.130 1542.740 448.450 ;
        RECT 1419.260 446.605 1419.400 448.130 ;
        RECT 1419.190 446.235 1419.470 446.605 ;
      LAYER via2 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
        RECT 1419.190 446.280 1419.470 446.560 ;
      LAYER met3 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
        RECT 1419.165 446.570 1419.495 446.585 ;
        RECT 1408.060 446.480 1419.495 446.570 ;
        RECT 1404.305 446.270 1419.495 446.480 ;
        RECT 1404.305 445.880 1408.305 446.270 ;
        RECT 1419.165 446.255 1419.495 446.270 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 1539.080 20.630 1539.140 ;
        RECT 113.690 1539.080 114.010 1539.140 ;
        RECT 20.310 1538.940 114.010 1539.080 ;
        RECT 20.310 1538.880 20.630 1538.940 ;
        RECT 113.690 1538.880 114.010 1538.940 ;
        RECT 113.690 1349.020 114.010 1349.080 ;
        RECT 383.710 1349.020 384.030 1349.080 ;
        RECT 113.690 1348.880 384.030 1349.020 ;
        RECT 113.690 1348.820 114.010 1348.880 ;
        RECT 383.710 1348.820 384.030 1348.880 ;
      LAYER via ;
        RECT 20.340 1538.880 20.600 1539.140 ;
        RECT 113.720 1538.880 113.980 1539.140 ;
        RECT 113.720 1348.820 113.980 1349.080 ;
        RECT 383.740 1348.820 384.000 1349.080 ;
      LAYER met2 ;
        RECT 20.330 1543.755 20.610 1544.125 ;
        RECT 20.400 1539.170 20.540 1543.755 ;
        RECT 20.340 1538.850 20.600 1539.170 ;
        RECT 113.720 1538.850 113.980 1539.170 ;
        RECT 113.780 1349.110 113.920 1538.850 ;
        RECT 113.720 1348.790 113.980 1349.110 ;
        RECT 383.740 1348.790 384.000 1349.110 ;
        RECT 383.800 1325.025 383.940 1348.790 ;
        RECT 383.690 1321.025 383.970 1325.025 ;
      LAYER via2 ;
        RECT 20.330 1543.800 20.610 1544.080 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 20.305 1544.090 20.635 1544.105 ;
        RECT -4.800 1543.790 20.635 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 20.305 1543.775 20.635 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 345.070 1340.860 345.390 1340.920 ;
        RECT 1416.410 1340.860 1416.730 1340.920 ;
        RECT 345.070 1340.720 1416.730 1340.860 ;
        RECT 345.070 1340.660 345.390 1340.720 ;
        RECT 1416.410 1340.660 1416.730 1340.720 ;
        RECT 19.390 1331.680 19.710 1331.740 ;
        RECT 345.070 1331.680 345.390 1331.740 ;
        RECT 19.390 1331.540 345.390 1331.680 ;
        RECT 19.390 1331.480 19.710 1331.540 ;
        RECT 345.070 1331.480 345.390 1331.540 ;
      LAYER via ;
        RECT 345.100 1340.660 345.360 1340.920 ;
        RECT 1416.440 1340.660 1416.700 1340.920 ;
        RECT 19.420 1331.480 19.680 1331.740 ;
        RECT 345.100 1331.480 345.360 1331.740 ;
      LAYER met2 ;
        RECT 345.100 1340.630 345.360 1340.950 ;
        RECT 1416.440 1340.630 1416.700 1340.950 ;
        RECT 345.160 1331.770 345.300 1340.630 ;
        RECT 19.420 1331.450 19.680 1331.770 ;
        RECT 345.100 1331.450 345.360 1331.770 ;
        RECT 19.480 1328.565 19.620 1331.450 ;
        RECT 19.410 1328.195 19.690 1328.565 ;
        RECT 1416.500 899.485 1416.640 1340.630 ;
        RECT 1416.430 899.115 1416.710 899.485 ;
      LAYER via2 ;
        RECT 19.410 1328.240 19.690 1328.520 ;
        RECT 1416.430 899.160 1416.710 899.440 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 19.385 1328.530 19.715 1328.545 ;
        RECT -4.800 1328.230 19.715 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 19.385 1328.215 19.715 1328.230 ;
        RECT 1416.405 899.450 1416.735 899.465 ;
        RECT 1408.060 899.360 1416.735 899.450 ;
        RECT 1404.305 899.150 1416.735 899.360 ;
        RECT 1404.305 898.760 1408.305 899.150 ;
        RECT 1416.405 899.135 1416.735 899.150 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 99.890 1339.840 100.210 1339.900 ;
        RECT 1145.470 1339.840 1145.790 1339.900 ;
        RECT 99.890 1339.700 1145.790 1339.840 ;
        RECT 99.890 1339.640 100.210 1339.700 ;
        RECT 1145.470 1339.640 1145.790 1339.700 ;
        RECT 14.790 1117.480 15.110 1117.540 ;
        RECT 99.890 1117.480 100.210 1117.540 ;
        RECT 14.790 1117.340 100.210 1117.480 ;
        RECT 14.790 1117.280 15.110 1117.340 ;
        RECT 99.890 1117.280 100.210 1117.340 ;
      LAYER via ;
        RECT 99.920 1339.640 100.180 1339.900 ;
        RECT 1145.500 1339.640 1145.760 1339.900 ;
        RECT 14.820 1117.280 15.080 1117.540 ;
        RECT 99.920 1117.280 100.180 1117.540 ;
      LAYER met2 ;
        RECT 99.920 1339.610 100.180 1339.930 ;
        RECT 1145.500 1339.610 1145.760 1339.930 ;
        RECT 99.980 1117.570 100.120 1339.610 ;
        RECT 1145.560 1325.025 1145.700 1339.610 ;
        RECT 1145.450 1321.025 1145.730 1325.025 ;
        RECT 14.820 1117.250 15.080 1117.570 ;
        RECT 99.920 1117.250 100.180 1117.570 ;
        RECT 14.880 1113.005 15.020 1117.250 ;
        RECT 14.810 1112.635 15.090 1113.005 ;
      LAYER via2 ;
        RECT 14.810 1112.680 15.090 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 14.785 1112.970 15.115 1112.985 ;
        RECT -4.800 1112.670 15.115 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 14.785 1112.655 15.115 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 903.195 20.610 903.565 ;
        RECT 20.400 897.445 20.540 903.195 ;
        RECT 20.330 897.075 20.610 897.445 ;
      LAYER via2 ;
        RECT 20.330 903.240 20.610 903.520 ;
        RECT 20.330 897.120 20.610 897.400 ;
      LAYER met3 ;
        RECT 1417.070 1107.220 1417.450 1107.540 ;
        RECT 1417.110 1106.180 1417.410 1107.220 ;
        RECT 1417.070 1105.860 1417.450 1106.180 ;
        RECT 1417.070 1046.020 1417.450 1046.340 ;
        RECT 1417.110 1044.980 1417.410 1046.020 ;
        RECT 1417.070 1044.660 1417.450 1044.980 ;
        RECT 20.305 903.530 20.635 903.545 ;
        RECT 306.630 903.530 307.010 903.540 ;
        RECT 20.305 903.230 307.010 903.530 ;
        RECT 20.305 903.215 20.635 903.230 ;
        RECT 306.630 903.220 307.010 903.230 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 20.305 897.410 20.635 897.425 ;
        RECT -4.800 897.110 20.635 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 20.305 897.095 20.635 897.110 ;
        RECT 1417.070 840.970 1417.450 840.980 ;
        RECT 1408.060 840.880 1417.450 840.970 ;
        RECT 1404.305 840.670 1417.450 840.880 ;
        RECT 1404.305 840.280 1408.305 840.670 ;
        RECT 1417.070 840.660 1417.450 840.670 ;
      LAYER via3 ;
        RECT 1417.100 1107.220 1417.420 1107.540 ;
        RECT 1417.100 1105.860 1417.420 1106.180 ;
        RECT 1417.100 1046.020 1417.420 1046.340 ;
        RECT 1417.100 1044.660 1417.420 1044.980 ;
        RECT 306.660 903.220 306.980 903.540 ;
        RECT 1417.100 840.660 1417.420 840.980 ;
      LAYER met4 ;
        RECT 306.230 1255.710 307.410 1256.890 ;
        RECT 1416.670 1255.710 1417.850 1256.890 ;
        RECT 306.670 903.545 306.970 1255.710 ;
        RECT 1417.110 1107.545 1417.410 1255.710 ;
        RECT 1417.095 1107.215 1417.425 1107.545 ;
        RECT 1417.095 1105.855 1417.425 1106.185 ;
        RECT 1417.110 1046.345 1417.410 1105.855 ;
        RECT 1417.095 1046.015 1417.425 1046.345 ;
        RECT 1417.095 1044.655 1417.425 1044.985 ;
        RECT 306.655 903.215 306.985 903.545 ;
        RECT 1417.110 840.985 1417.410 1044.655 ;
        RECT 1417.095 840.655 1417.425 840.985 ;
      LAYER met5 ;
        RECT 373.180 1265.700 416.180 1267.300 ;
        RECT 373.180 1257.100 374.780 1265.700 ;
        RECT 414.580 1260.500 416.180 1265.700 ;
        RECT 461.500 1265.700 502.660 1267.300 ;
        RECT 461.500 1263.900 463.100 1265.700 ;
        RECT 455.980 1262.300 463.100 1263.900 ;
        RECT 501.060 1263.900 502.660 1265.700 ;
        RECT 551.660 1265.700 563.380 1267.300 ;
        RECT 551.660 1263.900 553.260 1265.700 ;
        RECT 501.060 1262.300 510.940 1263.900 ;
        RECT 414.580 1258.900 425.380 1260.500 ;
        RECT 306.020 1255.500 374.780 1257.100 ;
        RECT 423.780 1257.100 425.380 1258.900 ;
        RECT 455.980 1257.100 457.580 1262.300 ;
        RECT 423.780 1255.500 457.580 1257.100 ;
        RECT 509.340 1260.500 510.940 1262.300 ;
        RECT 550.740 1262.300 553.260 1263.900 ;
        RECT 550.740 1260.500 552.340 1262.300 ;
        RECT 509.340 1258.900 552.340 1260.500 ;
        RECT 561.780 1260.500 563.380 1265.700 ;
        RECT 607.780 1265.700 654.460 1267.300 ;
        RECT 561.780 1258.900 604.780 1260.500 ;
        RECT 509.340 1255.500 511.860 1258.900 ;
        RECT 603.180 1257.100 604.780 1258.900 ;
        RECT 607.780 1257.100 609.380 1265.700 ;
        RECT 603.180 1255.500 609.380 1257.100 ;
        RECT 652.860 1257.100 654.460 1265.700 ;
        RECT 710.820 1265.700 776.820 1267.300 ;
        RECT 658.380 1258.900 701.380 1260.500 ;
        RECT 658.380 1257.100 659.980 1258.900 ;
        RECT 652.860 1255.500 659.980 1257.100 ;
        RECT 699.780 1257.100 701.380 1258.900 ;
        RECT 710.820 1257.100 712.420 1265.700 ;
        RECT 775.220 1260.500 776.820 1265.700 ;
        RECT 807.420 1265.700 873.420 1267.300 ;
        RECT 775.220 1258.900 798.900 1260.500 ;
        RECT 699.780 1255.500 712.420 1257.100 ;
        RECT 797.300 1257.100 798.900 1258.900 ;
        RECT 807.420 1257.100 809.020 1265.700 ;
        RECT 871.820 1260.500 873.420 1265.700 ;
        RECT 945.420 1265.700 993.020 1267.300 ;
        RECT 871.820 1258.900 895.500 1260.500 ;
        RECT 797.300 1255.500 809.020 1257.100 ;
        RECT 893.900 1257.100 895.500 1258.900 ;
        RECT 945.420 1257.100 947.020 1265.700 ;
        RECT 893.900 1255.500 922.180 1257.100 ;
        RECT 920.580 1253.700 922.180 1255.500 ;
        RECT 942.660 1255.500 947.020 1257.100 ;
        RECT 991.420 1257.100 993.020 1265.700 ;
        RECT 1049.380 1265.700 1096.060 1267.300 ;
        RECT 1049.380 1257.100 1050.980 1265.700 ;
        RECT 991.420 1255.500 1050.980 1257.100 ;
        RECT 1094.460 1257.100 1096.060 1265.700 ;
        RECT 1145.980 1265.700 1192.660 1267.300 ;
        RECT 1145.980 1257.100 1147.580 1265.700 ;
        RECT 1094.460 1255.500 1147.580 1257.100 ;
        RECT 1191.060 1257.100 1192.660 1265.700 ;
        RECT 1242.580 1265.700 1289.260 1267.300 ;
        RECT 1242.580 1257.100 1244.180 1265.700 ;
        RECT 1191.060 1255.500 1244.180 1257.100 ;
        RECT 1287.660 1257.100 1289.260 1265.700 ;
        RECT 1287.660 1255.500 1418.060 1257.100 ;
        RECT 942.660 1253.700 944.260 1255.500 ;
        RECT 920.580 1252.100 944.260 1253.700 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 19.850 676.500 20.170 676.560 ;
        RECT 265.490 676.500 265.810 676.560 ;
        RECT 19.850 676.360 265.810 676.500 ;
        RECT 19.850 676.300 20.170 676.360 ;
        RECT 265.490 676.300 265.810 676.360 ;
        RECT 265.490 212.740 265.810 212.800 ;
        RECT 732.390 212.740 732.710 212.800 ;
        RECT 265.490 212.600 732.710 212.740 ;
        RECT 265.490 212.540 265.810 212.600 ;
        RECT 732.390 212.540 732.710 212.600 ;
      LAYER via ;
        RECT 19.880 676.300 20.140 676.560 ;
        RECT 265.520 676.300 265.780 676.560 ;
        RECT 265.520 212.540 265.780 212.800 ;
        RECT 732.420 212.540 732.680 212.800 ;
      LAYER met2 ;
        RECT 19.870 681.515 20.150 681.885 ;
        RECT 19.940 676.590 20.080 681.515 ;
        RECT 19.880 676.270 20.140 676.590 ;
        RECT 265.520 676.270 265.780 676.590 ;
        RECT 265.580 212.830 265.720 676.270 ;
        RECT 732.370 216.000 732.650 220.000 ;
        RECT 732.480 212.830 732.620 216.000 ;
        RECT 265.520 212.510 265.780 212.830 ;
        RECT 732.420 212.510 732.680 212.830 ;
      LAYER via2 ;
        RECT 19.870 681.560 20.150 681.840 ;
      LAYER met3 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 19.845 681.850 20.175 681.865 ;
        RECT -4.800 681.550 20.175 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 19.845 681.535 20.175 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1404.305 1074.200 1408.305 1074.800 ;
        RECT 1407.910 1072.180 1408.210 1074.200 ;
        RECT 1407.870 1071.860 1408.250 1072.180 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 16.830 466.290 17.210 466.300 ;
        RECT -4.800 465.990 17.210 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 16.830 465.980 17.210 465.990 ;
        RECT 97.790 396.250 98.170 396.260 ;
        RECT 113.430 396.250 113.810 396.260 ;
        RECT 97.790 395.950 113.810 396.250 ;
        RECT 97.790 395.940 98.170 395.950 ;
        RECT 113.430 395.940 113.810 395.950 ;
        RECT 144.710 396.250 145.090 396.260 ;
        RECT 210.030 396.250 210.410 396.260 ;
        RECT 144.710 395.950 210.410 396.250 ;
        RECT 144.710 395.940 145.090 395.950 ;
        RECT 210.030 395.940 210.410 395.950 ;
      LAYER via3 ;
        RECT 1407.900 1071.860 1408.220 1072.180 ;
        RECT 16.860 465.980 17.180 466.300 ;
        RECT 97.820 395.940 98.140 396.260 ;
        RECT 113.460 395.940 113.780 396.260 ;
        RECT 144.740 395.940 145.060 396.260 ;
        RECT 210.060 395.940 210.380 396.260 ;
      LAYER met4 ;
        RECT 1407.895 1071.855 1408.225 1072.185 ;
        RECT 16.855 465.975 17.185 466.305 ;
        RECT 16.870 396.690 17.170 465.975 ;
        RECT 16.430 395.510 17.610 396.690 ;
        RECT 97.815 395.935 98.145 396.265 ;
        RECT 97.830 389.890 98.130 395.935 ;
        RECT 113.030 395.510 114.210 396.690 ;
        RECT 144.310 395.510 145.490 396.690 ;
        RECT 209.630 395.510 210.810 396.690 ;
        RECT 1407.910 396.250 1408.210 1071.855 ;
        RECT 1406.990 395.950 1408.210 396.250 ;
        RECT 1406.990 389.890 1407.290 395.950 ;
        RECT 97.390 388.710 98.570 389.890 ;
        RECT 1406.550 388.710 1407.730 389.890 ;
      LAYER met5 ;
        RECT 16.220 395.300 49.100 396.900 ;
        RECT 47.500 393.500 49.100 395.300 ;
        RECT 61.300 395.300 96.940 396.900 ;
        RECT 112.820 395.300 145.700 396.900 ;
        RECT 209.420 395.300 235.860 396.900 ;
        RECT 61.300 393.500 62.900 395.300 ;
        RECT 47.500 391.900 62.900 393.500 ;
        RECT 95.340 393.500 96.940 395.300 ;
        RECT 234.260 393.500 235.860 395.300 ;
        RECT 254.500 395.300 300.950 396.900 ;
        RECT 254.500 393.500 256.100 395.300 ;
        RECT 95.340 391.900 98.780 393.500 ;
        RECT 234.260 391.900 256.100 393.500 ;
        RECT 299.350 393.500 300.950 395.300 ;
        RECT 299.350 391.900 353.620 393.500 ;
        RECT 97.180 388.500 98.780 391.900 ;
        RECT 352.020 390.100 353.620 391.900 ;
        RECT 443.100 391.900 453.900 393.500 ;
        RECT 443.100 390.100 444.700 391.900 ;
        RECT 352.020 388.500 444.700 390.100 ;
        RECT 452.300 390.100 453.900 391.900 ;
        RECT 475.300 391.900 524.740 393.500 ;
        RECT 475.300 390.100 476.900 391.900 ;
        RECT 452.300 388.500 476.900 390.100 ;
        RECT 523.140 390.100 524.740 391.900 ;
        RECT 539.700 391.900 550.500 393.500 ;
        RECT 539.700 390.100 541.300 391.900 ;
        RECT 523.140 388.500 541.300 390.100 ;
        RECT 548.900 390.100 550.500 391.900 ;
        RECT 571.900 391.900 621.340 393.500 ;
        RECT 571.900 390.100 573.500 391.900 ;
        RECT 548.900 388.500 573.500 390.100 ;
        RECT 619.740 390.100 621.340 391.900 ;
        RECT 636.300 391.900 647.100 393.500 ;
        RECT 636.300 390.100 637.900 391.900 ;
        RECT 619.740 388.500 637.900 390.100 ;
        RECT 645.500 390.100 647.100 391.900 ;
        RECT 668.500 391.900 717.940 393.500 ;
        RECT 668.500 390.100 670.100 391.900 ;
        RECT 645.500 388.500 670.100 390.100 ;
        RECT 716.340 390.100 717.940 391.900 ;
        RECT 732.900 391.900 743.700 393.500 ;
        RECT 732.900 390.100 734.500 391.900 ;
        RECT 716.340 388.500 734.500 390.100 ;
        RECT 742.100 390.100 743.700 391.900 ;
        RECT 765.100 391.900 814.540 393.500 ;
        RECT 765.100 390.100 766.700 391.900 ;
        RECT 742.100 388.500 766.700 390.100 ;
        RECT 812.940 390.100 814.540 391.900 ;
        RECT 829.500 391.900 840.300 393.500 ;
        RECT 829.500 390.100 831.100 391.900 ;
        RECT 812.940 388.500 831.100 390.100 ;
        RECT 838.700 390.100 840.300 391.900 ;
        RECT 861.700 391.900 911.140 393.500 ;
        RECT 861.700 390.100 863.300 391.900 ;
        RECT 838.700 388.500 863.300 390.100 ;
        RECT 909.540 390.100 911.140 391.900 ;
        RECT 926.100 391.900 936.900 393.500 ;
        RECT 926.100 390.100 927.700 391.900 ;
        RECT 909.540 388.500 927.700 390.100 ;
        RECT 935.300 390.100 936.900 391.900 ;
        RECT 958.300 391.900 1007.740 393.500 ;
        RECT 958.300 390.100 959.900 391.900 ;
        RECT 935.300 388.500 959.900 390.100 ;
        RECT 1006.140 390.100 1007.740 391.900 ;
        RECT 1022.700 391.900 1033.500 393.500 ;
        RECT 1022.700 390.100 1024.300 391.900 ;
        RECT 1006.140 388.500 1024.300 390.100 ;
        RECT 1031.900 390.100 1033.500 391.900 ;
        RECT 1054.900 391.900 1104.340 393.500 ;
        RECT 1054.900 390.100 1056.500 391.900 ;
        RECT 1031.900 388.500 1056.500 390.100 ;
        RECT 1102.740 390.100 1104.340 391.900 ;
        RECT 1119.300 391.900 1130.100 393.500 ;
        RECT 1119.300 390.100 1120.900 391.900 ;
        RECT 1102.740 388.500 1120.900 390.100 ;
        RECT 1128.500 390.100 1130.100 391.900 ;
        RECT 1151.500 391.900 1200.940 393.500 ;
        RECT 1151.500 390.100 1153.100 391.900 ;
        RECT 1128.500 388.500 1153.100 390.100 ;
        RECT 1199.340 390.100 1200.940 391.900 ;
        RECT 1215.900 391.900 1226.700 393.500 ;
        RECT 1215.900 390.100 1217.500 391.900 ;
        RECT 1199.340 388.500 1217.500 390.100 ;
        RECT 1225.100 390.100 1226.700 391.900 ;
        RECT 1248.100 391.900 1297.540 393.500 ;
        RECT 1248.100 390.100 1249.700 391.900 ;
        RECT 1225.100 388.500 1249.700 390.100 ;
        RECT 1295.940 390.100 1297.540 391.900 ;
        RECT 1312.500 391.900 1323.300 393.500 ;
        RECT 1312.500 390.100 1314.100 391.900 ;
        RECT 1295.940 388.500 1314.100 390.100 ;
        RECT 1321.700 390.100 1323.300 391.900 ;
        RECT 1361.260 391.900 1407.940 393.500 ;
        RECT 1361.260 390.100 1362.860 391.900 ;
        RECT 1321.700 388.500 1362.860 390.100 ;
        RECT 1406.340 388.500 1407.940 391.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 210.360 17.870 210.420 ;
        RECT 444.890 210.360 445.210 210.420 ;
        RECT 17.550 210.220 445.210 210.360 ;
        RECT 17.550 210.160 17.870 210.220 ;
        RECT 444.890 210.160 445.210 210.220 ;
        RECT 444.890 206.280 445.210 206.340 ;
        RECT 485.830 206.280 486.150 206.340 ;
        RECT 444.890 206.140 486.150 206.280 ;
        RECT 444.890 206.080 445.210 206.140 ;
        RECT 485.830 206.080 486.150 206.140 ;
      LAYER via ;
        RECT 17.580 210.160 17.840 210.420 ;
        RECT 444.920 210.160 445.180 210.420 ;
        RECT 444.920 206.080 445.180 206.340 ;
        RECT 485.860 206.080 486.120 206.340 ;
      LAYER met2 ;
        RECT 17.570 250.395 17.850 250.765 ;
        RECT 17.640 210.450 17.780 250.395 ;
        RECT 485.810 216.000 486.090 220.000 ;
        RECT 17.580 210.130 17.840 210.450 ;
        RECT 444.920 210.130 445.180 210.450 ;
        RECT 444.980 206.370 445.120 210.130 ;
        RECT 485.920 206.370 486.060 216.000 ;
        RECT 444.920 206.050 445.180 206.370 ;
        RECT 485.860 206.050 486.120 206.370 ;
      LAYER via2 ;
        RECT 17.570 250.440 17.850 250.720 ;
      LAYER met3 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.545 250.730 17.875 250.745 ;
        RECT -4.800 250.430 17.875 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.545 250.415 17.875 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 30.890 517.720 31.210 517.780 ;
        RECT 296.770 517.720 297.090 517.780 ;
        RECT 30.890 517.580 297.090 517.720 ;
        RECT 30.890 517.520 31.210 517.580 ;
        RECT 296.770 517.520 297.090 517.580 ;
        RECT 14.790 36.960 15.110 37.020 ;
        RECT 30.890 36.960 31.210 37.020 ;
        RECT 14.790 36.820 31.210 36.960 ;
        RECT 14.790 36.760 15.110 36.820 ;
        RECT 30.890 36.760 31.210 36.820 ;
      LAYER via ;
        RECT 30.920 517.520 31.180 517.780 ;
        RECT 296.800 517.520 297.060 517.780 ;
        RECT 14.820 36.760 15.080 37.020 ;
        RECT 30.920 36.760 31.180 37.020 ;
      LAYER met2 ;
        RECT 296.790 519.675 297.070 520.045 ;
        RECT 296.860 517.810 297.000 519.675 ;
        RECT 30.920 517.490 31.180 517.810 ;
        RECT 296.800 517.490 297.060 517.810 ;
        RECT 30.980 37.050 31.120 517.490 ;
        RECT 14.820 36.730 15.080 37.050 ;
        RECT 30.920 36.730 31.180 37.050 ;
        RECT 14.880 35.885 15.020 36.730 ;
        RECT 14.810 35.515 15.090 35.885 ;
      LAYER via2 ;
        RECT 296.790 519.720 297.070 520.000 ;
        RECT 14.810 35.560 15.090 35.840 ;
      LAYER met3 ;
        RECT 296.765 520.010 297.095 520.025 ;
        RECT 296.765 519.920 310.500 520.010 ;
        RECT 296.765 519.710 314.000 519.920 ;
        RECT 296.765 519.695 297.095 519.710 ;
        RECT 310.000 519.320 314.000 519.710 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 14.785 35.850 15.115 35.865 ;
        RECT -4.800 35.550 15.115 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 14.785 35.535 15.115 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1057.150 1342.560 1057.470 1342.620 ;
        RECT 1466.550 1342.560 1466.870 1342.620 ;
        RECT 1057.150 1342.420 1466.870 1342.560 ;
        RECT 1057.150 1342.360 1057.470 1342.420 ;
        RECT 1466.550 1342.360 1466.870 1342.420 ;
        RECT 1466.550 910.760 1466.870 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 1466.550 910.620 2901.150 910.760 ;
        RECT 1466.550 910.560 1466.870 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 1057.180 1342.360 1057.440 1342.620 ;
        RECT 1466.580 1342.360 1466.840 1342.620 ;
        RECT 1466.580 910.560 1466.840 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 1057.180 1342.330 1057.440 1342.650 ;
        RECT 1466.580 1342.330 1466.840 1342.650 ;
        RECT 1057.240 1325.025 1057.380 1342.330 ;
        RECT 1057.130 1321.025 1057.410 1325.025 ;
        RECT 1466.640 910.850 1466.780 1342.330 ;
        RECT 1466.580 910.530 1466.840 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.770 210.360 642.090 210.420 ;
        RECT 2901.290 210.360 2901.610 210.420 ;
        RECT 641.770 210.220 2901.610 210.360 ;
        RECT 641.770 210.160 642.090 210.220 ;
        RECT 2901.290 210.160 2901.610 210.220 ;
        RECT 529.990 206.280 530.310 206.340 ;
        RECT 641.770 206.280 642.090 206.340 ;
        RECT 529.990 206.140 642.090 206.280 ;
        RECT 529.990 206.080 530.310 206.140 ;
        RECT 641.770 206.080 642.090 206.140 ;
      LAYER via ;
        RECT 641.800 210.160 642.060 210.420 ;
        RECT 2901.320 210.160 2901.580 210.420 ;
        RECT 530.020 206.080 530.280 206.340 ;
        RECT 641.800 206.080 642.060 206.340 ;
      LAYER met2 ;
        RECT 2901.310 1143.915 2901.590 1144.285 ;
        RECT 529.970 216.000 530.250 220.000 ;
        RECT 530.080 206.370 530.220 216.000 ;
        RECT 2901.380 210.450 2901.520 1143.915 ;
        RECT 641.800 210.130 642.060 210.450 ;
        RECT 2901.320 210.130 2901.580 210.450 ;
        RECT 641.860 206.370 642.000 210.130 ;
        RECT 530.020 206.050 530.280 206.370 ;
        RECT 641.800 206.050 642.060 206.370 ;
      LAYER via2 ;
        RECT 2901.310 1143.960 2901.590 1144.240 ;
      LAYER met3 ;
        RECT 2901.285 1144.250 2901.615 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2901.285 1143.950 2924.800 1144.250 ;
        RECT 2901.285 1143.935 2901.615 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1452.750 1373.500 1453.070 1373.560 ;
        RECT 2900.830 1373.500 2901.150 1373.560 ;
        RECT 1452.750 1373.360 2901.150 1373.500 ;
        RECT 1452.750 1373.300 1453.070 1373.360 ;
        RECT 2900.830 1373.300 2901.150 1373.360 ;
        RECT 925.590 213.080 925.910 213.140 ;
        RECT 1452.750 213.080 1453.070 213.140 ;
        RECT 925.590 212.940 1453.070 213.080 ;
        RECT 925.590 212.880 925.910 212.940 ;
        RECT 1452.750 212.880 1453.070 212.940 ;
      LAYER via ;
        RECT 1452.780 1373.300 1453.040 1373.560 ;
        RECT 2900.860 1373.300 2901.120 1373.560 ;
        RECT 925.620 212.880 925.880 213.140 ;
        RECT 1452.780 212.880 1453.040 213.140 ;
      LAYER met2 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
        RECT 2900.920 1373.590 2901.060 1378.515 ;
        RECT 1452.780 1373.270 1453.040 1373.590 ;
        RECT 2900.860 1373.270 2901.120 1373.590 ;
        RECT 925.570 216.000 925.850 220.000 ;
        RECT 925.680 213.170 925.820 216.000 ;
        RECT 1452.840 213.170 1452.980 1373.270 ;
        RECT 925.620 212.850 925.880 213.170 ;
        RECT 1452.780 212.850 1453.040 213.170 ;
      LAYER via2 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1459.650 1608.100 1459.970 1608.160 ;
        RECT 2900.830 1608.100 2901.150 1608.160 ;
        RECT 1459.650 1607.960 2901.150 1608.100 ;
        RECT 1459.650 1607.900 1459.970 1607.960 ;
        RECT 2900.830 1607.900 2901.150 1607.960 ;
        RECT 955.030 212.740 955.350 212.800 ;
        RECT 1459.650 212.740 1459.970 212.800 ;
        RECT 955.030 212.600 1459.970 212.740 ;
        RECT 955.030 212.540 955.350 212.600 ;
        RECT 1459.650 212.540 1459.970 212.600 ;
      LAYER via ;
        RECT 1459.680 1607.900 1459.940 1608.160 ;
        RECT 2900.860 1607.900 2901.120 1608.160 ;
        RECT 955.060 212.540 955.320 212.800 ;
        RECT 1459.680 212.540 1459.940 212.800 ;
      LAYER met2 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
        RECT 2900.920 1608.190 2901.060 1613.115 ;
        RECT 1459.680 1607.870 1459.940 1608.190 ;
        RECT 2900.860 1607.870 2901.120 1608.190 ;
        RECT 955.010 216.000 955.290 220.000 ;
        RECT 955.120 212.830 955.260 216.000 ;
        RECT 1459.740 212.830 1459.880 1607.870 ;
        RECT 955.060 212.510 955.320 212.830 ;
        RECT 1459.680 212.510 1459.940 212.830 ;
      LAYER via2 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
      LAYER met3 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 302.750 1842.700 303.070 1842.760 ;
        RECT 2900.830 1842.700 2901.150 1842.760 ;
        RECT 302.750 1842.560 2901.150 1842.700 ;
        RECT 302.750 1842.500 303.070 1842.560 ;
        RECT 2900.830 1842.500 2901.150 1842.560 ;
      LAYER via ;
        RECT 302.780 1842.500 303.040 1842.760 ;
        RECT 2900.860 1842.500 2901.120 1842.760 ;
      LAYER met2 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
        RECT 2900.920 1842.790 2901.060 1847.715 ;
        RECT 302.780 1842.470 303.040 1842.790 ;
        RECT 2900.860 1842.470 2901.120 1842.790 ;
        RECT 302.840 747.165 302.980 1842.470 ;
        RECT 302.770 746.795 303.050 747.165 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
        RECT 302.770 746.840 303.050 747.120 ;
      LAYER met3 ;
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 302.745 747.130 303.075 747.145 ;
        RECT 302.745 747.040 310.500 747.130 ;
        RECT 302.745 746.830 314.000 747.040 ;
        RECT 302.745 746.815 303.075 746.830 ;
        RECT 310.000 746.440 314.000 746.830 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1576.490 2077.300 1576.810 2077.360 ;
        RECT 2900.830 2077.300 2901.150 2077.360 ;
        RECT 1576.490 2077.160 2901.150 2077.300 ;
        RECT 1576.490 2077.100 1576.810 2077.160 ;
        RECT 2900.830 2077.100 2901.150 2077.160 ;
        RECT 1419.170 751.980 1419.490 752.040 ;
        RECT 1576.490 751.980 1576.810 752.040 ;
        RECT 1419.170 751.840 1576.810 751.980 ;
        RECT 1419.170 751.780 1419.490 751.840 ;
        RECT 1576.490 751.780 1576.810 751.840 ;
      LAYER via ;
        RECT 1576.520 2077.100 1576.780 2077.360 ;
        RECT 2900.860 2077.100 2901.120 2077.360 ;
        RECT 1419.200 751.780 1419.460 752.040 ;
        RECT 1576.520 751.780 1576.780 752.040 ;
      LAYER met2 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
        RECT 2900.920 2077.390 2901.060 2082.315 ;
        RECT 1576.520 2077.070 1576.780 2077.390 ;
        RECT 2900.860 2077.070 2901.120 2077.390 ;
        RECT 1576.580 752.070 1576.720 2077.070 ;
        RECT 1419.200 751.750 1419.460 752.070 ;
        RECT 1576.520 751.750 1576.780 752.070 ;
        RECT 1419.260 747.165 1419.400 751.750 ;
        RECT 1419.190 746.795 1419.470 747.165 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
        RECT 1419.190 746.840 1419.470 747.120 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 1419.165 747.130 1419.495 747.145 ;
        RECT 1408.060 747.040 1419.495 747.130 ;
        RECT 1404.305 746.830 1419.495 747.040 ;
        RECT 1404.305 746.440 1408.305 746.830 ;
        RECT 1419.165 746.815 1419.495 746.830 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 800.010 2311.900 800.330 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 800.010 2311.760 2901.150 2311.900 ;
        RECT 800.010 2311.700 800.330 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
        RECT 794.950 1332.020 795.270 1332.080 ;
        RECT 800.010 1332.020 800.330 1332.080 ;
        RECT 794.950 1331.880 800.330 1332.020 ;
        RECT 794.950 1331.820 795.270 1331.880 ;
        RECT 800.010 1331.820 800.330 1331.880 ;
      LAYER via ;
        RECT 800.040 2311.700 800.300 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
        RECT 794.980 1331.820 795.240 1332.080 ;
        RECT 800.040 1331.820 800.300 1332.080 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 800.040 2311.670 800.300 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 800.100 1332.110 800.240 2311.670 ;
        RECT 794.980 1331.790 795.240 1332.110 ;
        RECT 800.040 1331.790 800.300 1332.110 ;
        RECT 795.040 1325.025 795.180 1331.790 ;
        RECT 794.930 1321.025 795.210 1325.025 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 323.910 162.420 324.230 162.480 ;
        RECT 1116.030 162.420 1116.350 162.480 ;
        RECT 323.910 162.280 1116.350 162.420 ;
        RECT 323.910 162.220 324.230 162.280 ;
        RECT 1116.030 162.220 1116.350 162.280 ;
        RECT 1116.030 151.540 1116.350 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 1116.030 151.400 2901.150 151.540 ;
        RECT 1116.030 151.340 1116.350 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 323.940 162.220 324.200 162.480 ;
        RECT 1116.060 162.220 1116.320 162.480 ;
        RECT 1116.060 151.340 1116.320 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 322.050 216.650 322.330 220.000 ;
        RECT 322.050 216.510 324.140 216.650 ;
        RECT 322.050 216.000 322.330 216.510 ;
        RECT 324.000 162.510 324.140 216.510 ;
        RECT 323.940 162.190 324.200 162.510 ;
        RECT 1116.060 162.190 1116.320 162.510 ;
        RECT 1116.120 151.630 1116.260 162.190 ;
        RECT 1116.060 151.310 1116.320 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1472.990 2491.080 1473.310 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 1472.990 2490.940 2901.150 2491.080 ;
        RECT 1472.990 2490.880 1473.310 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
      LAYER via ;
        RECT 1473.020 2490.880 1473.280 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 1473.020 2490.850 1473.280 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 396.570 216.000 396.850 220.000 ;
        RECT 396.680 214.045 396.820 216.000 ;
        RECT 1473.080 214.045 1473.220 2490.850 ;
        RECT 396.610 213.675 396.890 214.045 ;
        RECT 1473.010 213.675 1473.290 214.045 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
        RECT 396.610 213.720 396.890 214.000 ;
        RECT 1473.010 213.720 1473.290 214.000 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 396.585 214.010 396.915 214.025 ;
        RECT 1472.985 214.010 1473.315 214.025 ;
        RECT 396.585 213.710 1473.315 214.010 ;
        RECT 396.585 213.695 396.915 213.710 ;
        RECT 1472.985 213.695 1473.315 213.710 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1407.210 2725.680 1407.530 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 1407.210 2725.540 2901.150 2725.680 ;
        RECT 1407.210 2725.480 1407.530 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
        RECT 1403.070 1338.480 1403.390 1338.540 ;
        RECT 1407.210 1338.480 1407.530 1338.540 ;
        RECT 1403.070 1338.340 1407.530 1338.480 ;
        RECT 1403.070 1338.280 1403.390 1338.340 ;
        RECT 1407.210 1338.280 1407.530 1338.340 ;
      LAYER via ;
        RECT 1407.240 2725.480 1407.500 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
        RECT 1403.100 1338.280 1403.360 1338.540 ;
        RECT 1407.240 1338.280 1407.500 1338.540 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 1407.240 2725.450 1407.500 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 1407.300 1338.570 1407.440 2725.450 ;
        RECT 1403.100 1338.250 1403.360 1338.570 ;
        RECT 1407.240 1338.250 1407.500 1338.570 ;
        RECT 1403.160 1325.025 1403.300 1338.250 ;
        RECT 1403.050 1321.025 1403.330 1325.025 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 365.310 2960.280 365.630 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 365.310 2960.140 2901.150 2960.280 ;
        RECT 365.310 2960.080 365.630 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 365.340 2960.080 365.600 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 365.340 2960.050 365.600 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 365.400 1325.050 365.540 2960.050 ;
        RECT 364.550 1325.025 365.540 1325.050 ;
        RECT 364.370 1324.910 365.540 1325.025 ;
        RECT 364.370 1321.025 364.650 1324.910 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1466.090 3194.880 1466.410 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 1466.090 3194.740 2901.150 3194.880 ;
        RECT 1466.090 3194.680 1466.410 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 1466.120 3194.680 1466.380 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 1466.120 3194.650 1466.380 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 806.890 216.000 807.170 220.000 ;
        RECT 807.000 212.005 807.140 216.000 ;
        RECT 1466.180 212.005 1466.320 3194.650 ;
        RECT 806.930 211.635 807.210 212.005 ;
        RECT 1466.110 211.635 1466.390 212.005 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
        RECT 806.930 211.680 807.210 211.960 ;
        RECT 1466.110 211.680 1466.390 211.960 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 806.905 211.970 807.235 211.985 ;
        RECT 1466.085 211.970 1466.415 211.985 ;
        RECT 806.905 211.670 1466.415 211.970 ;
        RECT 806.905 211.655 807.235 211.670 ;
        RECT 1466.085 211.655 1466.415 211.670 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1497.460 3429.680 1506.340 3429.820 ;
        RECT 1479.890 3429.480 1480.210 3429.540 ;
        RECT 1497.460 3429.480 1497.600 3429.680 ;
        RECT 1479.890 3429.340 1497.600 3429.480 ;
        RECT 1506.200 3429.480 1506.340 3429.680 ;
        RECT 2146.060 3429.680 2149.880 3429.820 ;
        RECT 2146.060 3429.480 2146.200 3429.680 ;
        RECT 1506.200 3429.340 2146.200 3429.480 ;
        RECT 2149.740 3429.480 2149.880 3429.680 ;
        RECT 2704.960 3429.680 2714.300 3429.820 ;
        RECT 2704.960 3429.480 2705.100 3429.680 ;
        RECT 2149.740 3429.340 2705.100 3429.480 ;
        RECT 2714.160 3429.480 2714.300 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2714.160 3429.340 2901.150 3429.480 ;
        RECT 1479.890 3429.280 1480.210 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
        RECT 411.310 199.140 411.630 199.200 ;
        RECT 1479.890 199.140 1480.210 199.200 ;
        RECT 411.310 199.000 1480.210 199.140 ;
        RECT 411.310 198.940 411.630 199.000 ;
        RECT 1479.890 198.940 1480.210 199.000 ;
      LAYER via ;
        RECT 1479.920 3429.280 1480.180 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
        RECT 411.340 198.940 411.600 199.200 ;
        RECT 1479.920 198.940 1480.180 199.200 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1479.920 3429.250 1480.180 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 411.290 216.000 411.570 220.000 ;
        RECT 411.400 199.230 411.540 216.000 ;
        RECT 1479.980 199.230 1480.120 3429.250 ;
        RECT 411.340 198.910 411.600 199.230 ;
        RECT 1479.920 198.910 1480.180 199.230 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2713.685 3332.765 2713.855 3422.355 ;
        RECT 2712.765 3008.405 2712.935 3042.915 ;
        RECT 2713.685 2946.525 2713.855 2994.635 ;
        RECT 2712.305 2753.065 2712.475 2801.175 ;
        RECT 2712.765 2428.705 2712.935 2463.215 ;
        RECT 2712.765 2331.805 2712.935 2366.655 ;
        RECT 2712.305 1993.845 2712.475 2028.355 ;
        RECT 2713.685 1766.725 2713.855 1787.635 ;
        RECT 2714.145 1703.825 2714.315 1766.215 ;
        RECT 2712.305 1400.885 2712.475 1448.995 ;
        RECT 2713.225 496.485 2713.395 507.195 ;
      LAYER mcon ;
        RECT 2713.685 3422.185 2713.855 3422.355 ;
        RECT 2712.765 3042.745 2712.935 3042.915 ;
        RECT 2713.685 2994.465 2713.855 2994.635 ;
        RECT 2712.305 2801.005 2712.475 2801.175 ;
        RECT 2712.765 2463.045 2712.935 2463.215 ;
        RECT 2712.765 2366.485 2712.935 2366.655 ;
        RECT 2712.305 2028.185 2712.475 2028.355 ;
        RECT 2713.685 1787.465 2713.855 1787.635 ;
        RECT 2714.145 1766.045 2714.315 1766.215 ;
        RECT 2712.305 1448.825 2712.475 1448.995 ;
        RECT 2713.225 507.025 2713.395 507.195 ;
      LAYER met1 ;
        RECT 2713.610 3491.360 2713.930 3491.420 ;
        RECT 2717.750 3491.360 2718.070 3491.420 ;
        RECT 2713.610 3491.220 2718.070 3491.360 ;
        RECT 2713.610 3491.160 2713.930 3491.220 ;
        RECT 2717.750 3491.160 2718.070 3491.220 ;
        RECT 2713.610 3443.220 2713.930 3443.480 ;
        RECT 2712.690 3443.080 2713.010 3443.140 ;
        RECT 2713.700 3443.080 2713.840 3443.220 ;
        RECT 2712.690 3442.940 2713.840 3443.080 ;
        RECT 2712.690 3442.880 2713.010 3442.940 ;
        RECT 2712.230 3422.340 2712.550 3422.400 ;
        RECT 2713.625 3422.340 2713.915 3422.385 ;
        RECT 2712.230 3422.200 2713.915 3422.340 ;
        RECT 2712.230 3422.140 2712.550 3422.200 ;
        RECT 2713.625 3422.155 2713.915 3422.200 ;
        RECT 2713.625 3332.920 2713.915 3332.965 ;
        RECT 2714.070 3332.920 2714.390 3332.980 ;
        RECT 2713.625 3332.780 2714.390 3332.920 ;
        RECT 2713.625 3332.735 2713.915 3332.780 ;
        RECT 2714.070 3332.720 2714.390 3332.780 ;
        RECT 2712.690 3236.360 2713.010 3236.420 ;
        RECT 2713.150 3236.360 2713.470 3236.420 ;
        RECT 2712.690 3236.220 2713.470 3236.360 ;
        RECT 2712.690 3236.160 2713.010 3236.220 ;
        RECT 2713.150 3236.160 2713.470 3236.220 ;
        RECT 2712.690 3202.020 2713.010 3202.080 ;
        RECT 2713.150 3202.020 2713.470 3202.080 ;
        RECT 2712.690 3201.880 2713.470 3202.020 ;
        RECT 2712.690 3201.820 2713.010 3201.880 ;
        RECT 2713.150 3201.820 2713.470 3201.880 ;
        RECT 2712.230 3153.400 2712.550 3153.460 ;
        RECT 2713.150 3153.400 2713.470 3153.460 ;
        RECT 2712.230 3153.260 2713.470 3153.400 ;
        RECT 2712.230 3153.200 2712.550 3153.260 ;
        RECT 2713.150 3153.200 2713.470 3153.260 ;
        RECT 2712.230 3056.840 2712.550 3056.900 ;
        RECT 2713.150 3056.840 2713.470 3056.900 ;
        RECT 2712.230 3056.700 2713.470 3056.840 ;
        RECT 2712.230 3056.640 2712.550 3056.700 ;
        RECT 2713.150 3056.640 2713.470 3056.700 ;
        RECT 2712.690 3042.900 2713.010 3042.960 ;
        RECT 2712.495 3042.760 2713.010 3042.900 ;
        RECT 2712.690 3042.700 2713.010 3042.760 ;
        RECT 2712.705 3008.560 2712.995 3008.605 ;
        RECT 2713.610 3008.560 2713.930 3008.620 ;
        RECT 2712.705 3008.420 2713.930 3008.560 ;
        RECT 2712.705 3008.375 2712.995 3008.420 ;
        RECT 2713.610 3008.360 2713.930 3008.420 ;
        RECT 2713.610 2994.620 2713.930 2994.680 ;
        RECT 2713.415 2994.480 2713.930 2994.620 ;
        RECT 2713.610 2994.420 2713.930 2994.480 ;
        RECT 2713.625 2946.680 2713.915 2946.725 ;
        RECT 2714.070 2946.680 2714.390 2946.740 ;
        RECT 2713.625 2946.540 2714.390 2946.680 ;
        RECT 2713.625 2946.495 2713.915 2946.540 ;
        RECT 2714.070 2946.480 2714.390 2946.540 ;
        RECT 2714.070 2912.340 2714.390 2912.400 ;
        RECT 2713.700 2912.200 2714.390 2912.340 ;
        RECT 2713.700 2911.720 2713.840 2912.200 ;
        RECT 2714.070 2912.140 2714.390 2912.200 ;
        RECT 2713.610 2911.460 2713.930 2911.720 ;
        RECT 2712.230 2815.580 2712.550 2815.840 ;
        RECT 2712.320 2815.160 2712.460 2815.580 ;
        RECT 2712.230 2814.900 2712.550 2815.160 ;
        RECT 2712.230 2801.160 2712.550 2801.220 ;
        RECT 2712.035 2801.020 2712.550 2801.160 ;
        RECT 2712.230 2800.960 2712.550 2801.020 ;
        RECT 2712.245 2753.220 2712.535 2753.265 ;
        RECT 2713.150 2753.220 2713.470 2753.280 ;
        RECT 2712.245 2753.080 2713.470 2753.220 ;
        RECT 2712.245 2753.035 2712.535 2753.080 ;
        RECT 2713.150 2753.020 2713.470 2753.080 ;
        RECT 2712.230 2718.200 2712.550 2718.260 ;
        RECT 2713.150 2718.200 2713.470 2718.260 ;
        RECT 2712.230 2718.060 2713.470 2718.200 ;
        RECT 2712.230 2718.000 2712.550 2718.060 ;
        RECT 2713.150 2718.000 2713.470 2718.060 ;
        RECT 2712.230 2670.260 2712.550 2670.320 ;
        RECT 2713.150 2670.260 2713.470 2670.320 ;
        RECT 2712.230 2670.120 2713.470 2670.260 ;
        RECT 2712.230 2670.060 2712.550 2670.120 ;
        RECT 2713.150 2670.060 2713.470 2670.120 ;
        RECT 2713.150 2622.120 2713.470 2622.380 ;
        RECT 2713.240 2621.980 2713.380 2622.120 ;
        RECT 2713.610 2621.980 2713.930 2622.040 ;
        RECT 2713.240 2621.840 2713.930 2621.980 ;
        RECT 2713.610 2621.780 2713.930 2621.840 ;
        RECT 2712.690 2560.100 2713.010 2560.160 ;
        RECT 2714.070 2560.100 2714.390 2560.160 ;
        RECT 2712.690 2559.960 2714.390 2560.100 ;
        RECT 2712.690 2559.900 2713.010 2559.960 ;
        RECT 2714.070 2559.900 2714.390 2559.960 ;
        RECT 2713.150 2511.820 2713.470 2511.880 ;
        RECT 2714.070 2511.820 2714.390 2511.880 ;
        RECT 2713.150 2511.680 2714.390 2511.820 ;
        RECT 2713.150 2511.620 2713.470 2511.680 ;
        RECT 2714.070 2511.620 2714.390 2511.680 ;
        RECT 2712.690 2463.200 2713.010 2463.260 ;
        RECT 2712.495 2463.060 2713.010 2463.200 ;
        RECT 2712.690 2463.000 2713.010 2463.060 ;
        RECT 2712.690 2428.860 2713.010 2428.920 ;
        RECT 2712.495 2428.720 2713.010 2428.860 ;
        RECT 2712.690 2428.660 2713.010 2428.720 ;
        RECT 2712.230 2380.580 2712.550 2380.640 ;
        RECT 2713.150 2380.580 2713.470 2380.640 ;
        RECT 2712.230 2380.440 2713.470 2380.580 ;
        RECT 2712.230 2380.380 2712.550 2380.440 ;
        RECT 2713.150 2380.380 2713.470 2380.440 ;
        RECT 2712.690 2366.640 2713.010 2366.700 ;
        RECT 2712.495 2366.500 2713.010 2366.640 ;
        RECT 2712.690 2366.440 2713.010 2366.500 ;
        RECT 2712.690 2331.960 2713.010 2332.020 ;
        RECT 2712.495 2331.820 2713.010 2331.960 ;
        RECT 2712.690 2331.760 2713.010 2331.820 ;
        RECT 2711.770 2235.540 2712.090 2235.800 ;
        RECT 2711.860 2235.400 2712.000 2235.540 ;
        RECT 2712.230 2235.400 2712.550 2235.460 ;
        RECT 2711.860 2235.260 2712.550 2235.400 ;
        RECT 2712.230 2235.200 2712.550 2235.260 ;
        RECT 2710.850 2221.800 2711.170 2221.860 ;
        RECT 2712.230 2221.800 2712.550 2221.860 ;
        RECT 2710.850 2221.660 2712.550 2221.800 ;
        RECT 2710.850 2221.600 2711.170 2221.660 ;
        RECT 2712.230 2221.600 2712.550 2221.660 ;
        RECT 2711.770 2138.980 2712.090 2139.240 ;
        RECT 2711.860 2138.840 2712.000 2138.980 ;
        RECT 2712.230 2138.840 2712.550 2138.900 ;
        RECT 2711.860 2138.700 2712.550 2138.840 ;
        RECT 2712.230 2138.640 2712.550 2138.700 ;
        RECT 2710.850 2125.240 2711.170 2125.300 ;
        RECT 2712.230 2125.240 2712.550 2125.300 ;
        RECT 2710.850 2125.100 2712.550 2125.240 ;
        RECT 2710.850 2125.040 2711.170 2125.100 ;
        RECT 2712.230 2125.040 2712.550 2125.100 ;
        RECT 2711.770 2042.420 2712.090 2042.680 ;
        RECT 2711.860 2041.940 2712.000 2042.420 ;
        RECT 2712.230 2041.940 2712.550 2042.000 ;
        RECT 2711.860 2041.800 2712.550 2041.940 ;
        RECT 2712.230 2041.740 2712.550 2041.800 ;
        RECT 2712.230 2028.340 2712.550 2028.400 ;
        RECT 2712.035 2028.200 2712.550 2028.340 ;
        RECT 2712.230 2028.140 2712.550 2028.200 ;
        RECT 2712.230 1994.000 2712.550 1994.060 ;
        RECT 2712.035 1993.860 2712.550 1994.000 ;
        RECT 2712.230 1993.800 2712.550 1993.860 ;
        RECT 2712.230 1945.860 2712.550 1946.120 ;
        RECT 2712.320 1945.440 2712.460 1945.860 ;
        RECT 2712.230 1945.180 2712.550 1945.440 ;
        RECT 2712.230 1897.440 2712.550 1897.500 ;
        RECT 2713.150 1897.440 2713.470 1897.500 ;
        RECT 2712.230 1897.300 2713.470 1897.440 ;
        RECT 2712.230 1897.240 2712.550 1897.300 ;
        RECT 2713.150 1897.240 2713.470 1897.300 ;
        RECT 2713.610 1787.620 2713.930 1787.680 ;
        RECT 2713.415 1787.480 2713.930 1787.620 ;
        RECT 2713.610 1787.420 2713.930 1787.480 ;
        RECT 2713.610 1766.880 2713.930 1766.940 ;
        RECT 2713.415 1766.740 2713.930 1766.880 ;
        RECT 2713.610 1766.680 2713.930 1766.740 ;
        RECT 2714.070 1766.200 2714.390 1766.260 ;
        RECT 2713.875 1766.060 2714.390 1766.200 ;
        RECT 2714.070 1766.000 2714.390 1766.060 ;
        RECT 2714.070 1703.980 2714.390 1704.040 ;
        RECT 2713.875 1703.840 2714.390 1703.980 ;
        RECT 2714.070 1703.780 2714.390 1703.840 ;
        RECT 2713.150 1628.500 2713.470 1628.560 ;
        RECT 2713.610 1628.500 2713.930 1628.560 ;
        RECT 2713.150 1628.360 2713.930 1628.500 ;
        RECT 2713.150 1628.300 2713.470 1628.360 ;
        RECT 2713.610 1628.300 2713.930 1628.360 ;
        RECT 2712.690 1594.160 2713.010 1594.220 ;
        RECT 2713.150 1594.160 2713.470 1594.220 ;
        RECT 2712.690 1594.020 2713.470 1594.160 ;
        RECT 2712.690 1593.960 2713.010 1594.020 ;
        RECT 2713.150 1593.960 2713.470 1594.020 ;
        RECT 2712.690 1559.820 2713.010 1559.880 ;
        RECT 2713.150 1559.820 2713.470 1559.880 ;
        RECT 2712.690 1559.680 2713.470 1559.820 ;
        RECT 2712.690 1559.620 2713.010 1559.680 ;
        RECT 2713.150 1559.620 2713.470 1559.680 ;
        RECT 2712.230 1511.200 2712.550 1511.260 ;
        RECT 2713.150 1511.200 2713.470 1511.260 ;
        RECT 2712.230 1511.060 2713.470 1511.200 ;
        RECT 2712.230 1511.000 2712.550 1511.060 ;
        RECT 2713.150 1511.000 2713.470 1511.060 ;
        RECT 2712.245 1448.980 2712.535 1449.025 ;
        RECT 2713.150 1448.980 2713.470 1449.040 ;
        RECT 2712.245 1448.840 2713.470 1448.980 ;
        RECT 2712.245 1448.795 2712.535 1448.840 ;
        RECT 2713.150 1448.780 2713.470 1448.840 ;
        RECT 2712.230 1401.040 2712.550 1401.100 ;
        RECT 2712.035 1400.900 2712.550 1401.040 ;
        RECT 2712.230 1400.840 2712.550 1400.900 ;
        RECT 2711.770 1338.820 2712.090 1338.880 ;
        RECT 2713.150 1338.820 2713.470 1338.880 ;
        RECT 2711.770 1338.680 2713.470 1338.820 ;
        RECT 2711.770 1338.620 2712.090 1338.680 ;
        RECT 2713.150 1338.620 2713.470 1338.680 ;
        RECT 2711.770 1221.180 2712.090 1221.240 ;
        RECT 2713.150 1221.180 2713.470 1221.240 ;
        RECT 2711.770 1221.040 2713.470 1221.180 ;
        RECT 2711.770 1220.980 2712.090 1221.040 ;
        RECT 2713.150 1220.980 2713.470 1221.040 ;
        RECT 2712.690 1159.300 2713.010 1159.360 ;
        RECT 2713.610 1159.300 2713.930 1159.360 ;
        RECT 2712.690 1159.160 2713.930 1159.300 ;
        RECT 2712.690 1159.100 2713.010 1159.160 ;
        RECT 2713.610 1159.100 2713.930 1159.160 ;
        RECT 2711.770 1111.020 2712.090 1111.080 ;
        RECT 2713.150 1111.020 2713.470 1111.080 ;
        RECT 2711.770 1110.880 2713.470 1111.020 ;
        RECT 2711.770 1110.820 2712.090 1110.880 ;
        RECT 2713.150 1110.820 2713.470 1110.880 ;
        RECT 2712.690 1014.460 2713.010 1014.520 ;
        RECT 2713.150 1014.460 2713.470 1014.520 ;
        RECT 2712.690 1014.320 2713.470 1014.460 ;
        RECT 2712.690 1014.260 2713.010 1014.320 ;
        RECT 2713.150 1014.260 2713.470 1014.320 ;
        RECT 2713.150 979.920 2713.470 980.180 ;
        RECT 2713.240 979.780 2713.380 979.920 ;
        RECT 2713.610 979.780 2713.930 979.840 ;
        RECT 2713.240 979.640 2713.930 979.780 ;
        RECT 2713.610 979.580 2713.930 979.640 ;
        RECT 2712.690 917.900 2713.010 917.960 ;
        RECT 2714.070 917.900 2714.390 917.960 ;
        RECT 2712.690 917.760 2714.390 917.900 ;
        RECT 2712.690 917.700 2713.010 917.760 ;
        RECT 2714.070 917.700 2714.390 917.760 ;
        RECT 2713.150 869.620 2713.470 869.680 ;
        RECT 2714.070 869.620 2714.390 869.680 ;
        RECT 2713.150 869.480 2714.390 869.620 ;
        RECT 2713.150 869.420 2713.470 869.480 ;
        RECT 2714.070 869.420 2714.390 869.480 ;
        RECT 2711.770 845.480 2712.090 845.540 ;
        RECT 2713.150 845.480 2713.470 845.540 ;
        RECT 2711.770 845.340 2713.470 845.480 ;
        RECT 2711.770 845.280 2712.090 845.340 ;
        RECT 2713.150 845.280 2713.470 845.340 ;
        RECT 2711.770 807.060 2712.090 807.120 ;
        RECT 2713.150 807.060 2713.470 807.120 ;
        RECT 2711.770 806.920 2713.470 807.060 ;
        RECT 2711.770 806.860 2712.090 806.920 ;
        RECT 2713.150 806.860 2713.470 806.920 ;
        RECT 2711.770 759.120 2712.090 759.180 ;
        RECT 2713.150 759.120 2713.470 759.180 ;
        RECT 2711.770 758.980 2713.470 759.120 ;
        RECT 2711.770 758.920 2712.090 758.980 ;
        RECT 2713.150 758.920 2713.470 758.980 ;
        RECT 2711.770 710.500 2712.090 710.560 ;
        RECT 2713.150 710.500 2713.470 710.560 ;
        RECT 2711.770 710.360 2713.470 710.500 ;
        RECT 2711.770 710.300 2712.090 710.360 ;
        RECT 2713.150 710.300 2713.470 710.360 ;
        RECT 2711.770 662.560 2712.090 662.620 ;
        RECT 2713.150 662.560 2713.470 662.620 ;
        RECT 2711.770 662.420 2713.470 662.560 ;
        RECT 2711.770 662.360 2712.090 662.420 ;
        RECT 2713.150 662.360 2713.470 662.420 ;
        RECT 2711.770 641.480 2712.090 641.540 ;
        RECT 2713.150 641.480 2713.470 641.540 ;
        RECT 2711.770 641.340 2713.470 641.480 ;
        RECT 2711.770 641.280 2712.090 641.340 ;
        RECT 2713.150 641.280 2713.470 641.340 ;
        RECT 2711.770 579.600 2712.090 579.660 ;
        RECT 2712.690 579.600 2713.010 579.660 ;
        RECT 2711.770 579.460 2713.010 579.600 ;
        RECT 2711.770 579.400 2712.090 579.460 ;
        RECT 2712.690 579.400 2713.010 579.460 ;
        RECT 2713.150 507.180 2713.470 507.240 ;
        RECT 2712.955 507.040 2713.470 507.180 ;
        RECT 2713.150 506.980 2713.470 507.040 ;
        RECT 2713.165 496.640 2713.455 496.685 ;
        RECT 2713.610 496.640 2713.930 496.700 ;
        RECT 2713.165 496.500 2713.930 496.640 ;
        RECT 2713.165 496.455 2713.455 496.500 ;
        RECT 2713.610 496.440 2713.930 496.500 ;
        RECT 2712.690 337.860 2713.010 337.920 ;
        RECT 2713.610 337.860 2713.930 337.920 ;
        RECT 2712.690 337.720 2713.930 337.860 ;
        RECT 2712.690 337.660 2713.010 337.720 ;
        RECT 2713.610 337.660 2713.930 337.720 ;
        RECT 519.870 205.600 520.190 205.660 ;
        RECT 607.270 205.600 607.590 205.660 ;
        RECT 519.870 205.460 607.590 205.600 ;
        RECT 519.870 205.400 520.190 205.460 ;
        RECT 607.270 205.400 607.590 205.460 ;
      LAYER via ;
        RECT 2713.640 3491.160 2713.900 3491.420 ;
        RECT 2717.780 3491.160 2718.040 3491.420 ;
        RECT 2713.640 3443.220 2713.900 3443.480 ;
        RECT 2712.720 3442.880 2712.980 3443.140 ;
        RECT 2712.260 3422.140 2712.520 3422.400 ;
        RECT 2714.100 3332.720 2714.360 3332.980 ;
        RECT 2712.720 3236.160 2712.980 3236.420 ;
        RECT 2713.180 3236.160 2713.440 3236.420 ;
        RECT 2712.720 3201.820 2712.980 3202.080 ;
        RECT 2713.180 3201.820 2713.440 3202.080 ;
        RECT 2712.260 3153.200 2712.520 3153.460 ;
        RECT 2713.180 3153.200 2713.440 3153.460 ;
        RECT 2712.260 3056.640 2712.520 3056.900 ;
        RECT 2713.180 3056.640 2713.440 3056.900 ;
        RECT 2712.720 3042.700 2712.980 3042.960 ;
        RECT 2713.640 3008.360 2713.900 3008.620 ;
        RECT 2713.640 2994.420 2713.900 2994.680 ;
        RECT 2714.100 2946.480 2714.360 2946.740 ;
        RECT 2714.100 2912.140 2714.360 2912.400 ;
        RECT 2713.640 2911.460 2713.900 2911.720 ;
        RECT 2712.260 2815.580 2712.520 2815.840 ;
        RECT 2712.260 2814.900 2712.520 2815.160 ;
        RECT 2712.260 2800.960 2712.520 2801.220 ;
        RECT 2713.180 2753.020 2713.440 2753.280 ;
        RECT 2712.260 2718.000 2712.520 2718.260 ;
        RECT 2713.180 2718.000 2713.440 2718.260 ;
        RECT 2712.260 2670.060 2712.520 2670.320 ;
        RECT 2713.180 2670.060 2713.440 2670.320 ;
        RECT 2713.180 2622.120 2713.440 2622.380 ;
        RECT 2713.640 2621.780 2713.900 2622.040 ;
        RECT 2712.720 2559.900 2712.980 2560.160 ;
        RECT 2714.100 2559.900 2714.360 2560.160 ;
        RECT 2713.180 2511.620 2713.440 2511.880 ;
        RECT 2714.100 2511.620 2714.360 2511.880 ;
        RECT 2712.720 2463.000 2712.980 2463.260 ;
        RECT 2712.720 2428.660 2712.980 2428.920 ;
        RECT 2712.260 2380.380 2712.520 2380.640 ;
        RECT 2713.180 2380.380 2713.440 2380.640 ;
        RECT 2712.720 2366.440 2712.980 2366.700 ;
        RECT 2712.720 2331.760 2712.980 2332.020 ;
        RECT 2711.800 2235.540 2712.060 2235.800 ;
        RECT 2712.260 2235.200 2712.520 2235.460 ;
        RECT 2710.880 2221.600 2711.140 2221.860 ;
        RECT 2712.260 2221.600 2712.520 2221.860 ;
        RECT 2711.800 2138.980 2712.060 2139.240 ;
        RECT 2712.260 2138.640 2712.520 2138.900 ;
        RECT 2710.880 2125.040 2711.140 2125.300 ;
        RECT 2712.260 2125.040 2712.520 2125.300 ;
        RECT 2711.800 2042.420 2712.060 2042.680 ;
        RECT 2712.260 2041.740 2712.520 2042.000 ;
        RECT 2712.260 2028.140 2712.520 2028.400 ;
        RECT 2712.260 1993.800 2712.520 1994.060 ;
        RECT 2712.260 1945.860 2712.520 1946.120 ;
        RECT 2712.260 1945.180 2712.520 1945.440 ;
        RECT 2712.260 1897.240 2712.520 1897.500 ;
        RECT 2713.180 1897.240 2713.440 1897.500 ;
        RECT 2713.640 1787.420 2713.900 1787.680 ;
        RECT 2713.640 1766.680 2713.900 1766.940 ;
        RECT 2714.100 1766.000 2714.360 1766.260 ;
        RECT 2714.100 1703.780 2714.360 1704.040 ;
        RECT 2713.180 1628.300 2713.440 1628.560 ;
        RECT 2713.640 1628.300 2713.900 1628.560 ;
        RECT 2712.720 1593.960 2712.980 1594.220 ;
        RECT 2713.180 1593.960 2713.440 1594.220 ;
        RECT 2712.720 1559.620 2712.980 1559.880 ;
        RECT 2713.180 1559.620 2713.440 1559.880 ;
        RECT 2712.260 1511.000 2712.520 1511.260 ;
        RECT 2713.180 1511.000 2713.440 1511.260 ;
        RECT 2713.180 1448.780 2713.440 1449.040 ;
        RECT 2712.260 1400.840 2712.520 1401.100 ;
        RECT 2711.800 1338.620 2712.060 1338.880 ;
        RECT 2713.180 1338.620 2713.440 1338.880 ;
        RECT 2711.800 1220.980 2712.060 1221.240 ;
        RECT 2713.180 1220.980 2713.440 1221.240 ;
        RECT 2712.720 1159.100 2712.980 1159.360 ;
        RECT 2713.640 1159.100 2713.900 1159.360 ;
        RECT 2711.800 1110.820 2712.060 1111.080 ;
        RECT 2713.180 1110.820 2713.440 1111.080 ;
        RECT 2712.720 1014.260 2712.980 1014.520 ;
        RECT 2713.180 1014.260 2713.440 1014.520 ;
        RECT 2713.180 979.920 2713.440 980.180 ;
        RECT 2713.640 979.580 2713.900 979.840 ;
        RECT 2712.720 917.700 2712.980 917.960 ;
        RECT 2714.100 917.700 2714.360 917.960 ;
        RECT 2713.180 869.420 2713.440 869.680 ;
        RECT 2714.100 869.420 2714.360 869.680 ;
        RECT 2711.800 845.280 2712.060 845.540 ;
        RECT 2713.180 845.280 2713.440 845.540 ;
        RECT 2711.800 806.860 2712.060 807.120 ;
        RECT 2713.180 806.860 2713.440 807.120 ;
        RECT 2711.800 758.920 2712.060 759.180 ;
        RECT 2713.180 758.920 2713.440 759.180 ;
        RECT 2711.800 710.300 2712.060 710.560 ;
        RECT 2713.180 710.300 2713.440 710.560 ;
        RECT 2711.800 662.360 2712.060 662.620 ;
        RECT 2713.180 662.360 2713.440 662.620 ;
        RECT 2711.800 641.280 2712.060 641.540 ;
        RECT 2713.180 641.280 2713.440 641.540 ;
        RECT 2711.800 579.400 2712.060 579.660 ;
        RECT 2712.720 579.400 2712.980 579.660 ;
        RECT 2713.180 506.980 2713.440 507.240 ;
        RECT 2713.640 496.440 2713.900 496.700 ;
        RECT 2712.720 337.660 2712.980 337.920 ;
        RECT 2713.640 337.660 2713.900 337.920 ;
        RECT 519.900 205.400 520.160 205.660 ;
        RECT 607.300 205.400 607.560 205.660 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3517.370 2717.520 3517.600 ;
        RECT 2717.380 3517.230 2717.980 3517.370 ;
        RECT 2717.840 3491.450 2717.980 3517.230 ;
        RECT 2713.640 3491.130 2713.900 3491.450 ;
        RECT 2717.780 3491.130 2718.040 3491.450 ;
        RECT 2713.700 3443.510 2713.840 3491.130 ;
        RECT 2713.640 3443.190 2713.900 3443.510 ;
        RECT 2712.720 3442.850 2712.980 3443.170 ;
        RECT 2712.780 3429.650 2712.920 3442.850 ;
        RECT 2712.320 3429.510 2712.920 3429.650 ;
        RECT 2712.320 3422.430 2712.460 3429.510 ;
        RECT 2712.260 3422.110 2712.520 3422.430 ;
        RECT 2714.100 3332.690 2714.360 3333.010 ;
        RECT 2714.160 3298.410 2714.300 3332.690 ;
        RECT 2713.240 3298.270 2714.300 3298.410 ;
        RECT 2713.240 3236.450 2713.380 3298.270 ;
        RECT 2712.720 3236.130 2712.980 3236.450 ;
        RECT 2713.180 3236.130 2713.440 3236.450 ;
        RECT 2712.780 3202.110 2712.920 3236.130 ;
        RECT 2712.720 3201.790 2712.980 3202.110 ;
        RECT 2713.180 3201.790 2713.440 3202.110 ;
        RECT 2713.240 3153.490 2713.380 3201.790 ;
        RECT 2712.260 3153.170 2712.520 3153.490 ;
        RECT 2713.180 3153.170 2713.440 3153.490 ;
        RECT 2712.320 3152.890 2712.460 3153.170 ;
        RECT 2712.320 3152.750 2712.920 3152.890 ;
        RECT 2712.780 3105.290 2712.920 3152.750 ;
        RECT 2712.780 3105.150 2713.380 3105.290 ;
        RECT 2713.240 3056.930 2713.380 3105.150 ;
        RECT 2712.260 3056.610 2712.520 3056.930 ;
        RECT 2713.180 3056.610 2713.440 3056.930 ;
        RECT 2712.320 3056.330 2712.460 3056.610 ;
        RECT 2712.320 3056.190 2712.920 3056.330 ;
        RECT 2712.780 3042.990 2712.920 3056.190 ;
        RECT 2712.720 3042.670 2712.980 3042.990 ;
        RECT 2713.640 3008.330 2713.900 3008.650 ;
        RECT 2713.700 2994.710 2713.840 3008.330 ;
        RECT 2713.640 2994.390 2713.900 2994.710 ;
        RECT 2714.100 2946.450 2714.360 2946.770 ;
        RECT 2714.160 2912.430 2714.300 2946.450 ;
        RECT 2714.100 2912.110 2714.360 2912.430 ;
        RECT 2713.640 2911.430 2713.900 2911.750 ;
        RECT 2713.700 2863.210 2713.840 2911.430 ;
        RECT 2712.780 2863.070 2713.840 2863.210 ;
        RECT 2712.780 2849.610 2712.920 2863.070 ;
        RECT 2712.320 2849.470 2712.920 2849.610 ;
        RECT 2712.320 2815.870 2712.460 2849.470 ;
        RECT 2712.260 2815.550 2712.520 2815.870 ;
        RECT 2712.260 2814.870 2712.520 2815.190 ;
        RECT 2712.320 2801.250 2712.460 2814.870 ;
        RECT 2712.260 2800.930 2712.520 2801.250 ;
        RECT 2713.180 2752.990 2713.440 2753.310 ;
        RECT 2713.240 2718.290 2713.380 2752.990 ;
        RECT 2712.260 2717.970 2712.520 2718.290 ;
        RECT 2713.180 2717.970 2713.440 2718.290 ;
        RECT 2712.320 2670.350 2712.460 2717.970 ;
        RECT 2712.260 2670.030 2712.520 2670.350 ;
        RECT 2713.180 2670.030 2713.440 2670.350 ;
        RECT 2713.240 2622.410 2713.380 2670.030 ;
        RECT 2713.180 2622.090 2713.440 2622.410 ;
        RECT 2713.640 2621.750 2713.900 2622.070 ;
        RECT 2713.700 2608.325 2713.840 2621.750 ;
        RECT 2712.710 2607.955 2712.990 2608.325 ;
        RECT 2713.630 2607.955 2713.910 2608.325 ;
        RECT 2712.780 2560.190 2712.920 2607.955 ;
        RECT 2712.720 2559.870 2712.980 2560.190 ;
        RECT 2714.100 2559.870 2714.360 2560.190 ;
        RECT 2714.160 2511.910 2714.300 2559.870 ;
        RECT 2713.180 2511.765 2713.440 2511.910 ;
        RECT 2711.790 2511.395 2712.070 2511.765 ;
        RECT 2713.170 2511.395 2713.450 2511.765 ;
        RECT 2714.100 2511.590 2714.360 2511.910 ;
        RECT 2711.860 2463.485 2712.000 2511.395 ;
        RECT 2711.790 2463.115 2712.070 2463.485 ;
        RECT 2712.710 2463.115 2712.990 2463.485 ;
        RECT 2712.720 2462.970 2712.980 2463.115 ;
        RECT 2712.720 2428.630 2712.980 2428.950 ;
        RECT 2712.780 2415.090 2712.920 2428.630 ;
        RECT 2712.780 2414.950 2713.380 2415.090 ;
        RECT 2713.240 2380.670 2713.380 2414.950 ;
        RECT 2712.260 2380.410 2712.520 2380.670 ;
        RECT 2712.260 2380.350 2712.920 2380.410 ;
        RECT 2713.180 2380.350 2713.440 2380.670 ;
        RECT 2712.320 2380.270 2712.920 2380.350 ;
        RECT 2712.780 2366.730 2712.920 2380.270 ;
        RECT 2712.720 2366.410 2712.980 2366.730 ;
        RECT 2712.720 2331.730 2712.980 2332.050 ;
        RECT 2712.780 2318.530 2712.920 2331.730 ;
        RECT 2712.780 2318.390 2713.380 2318.530 ;
        RECT 2713.240 2270.365 2713.380 2318.390 ;
        RECT 2711.790 2269.995 2712.070 2270.365 ;
        RECT 2713.170 2269.995 2713.450 2270.365 ;
        RECT 2711.860 2235.830 2712.000 2269.995 ;
        RECT 2711.800 2235.510 2712.060 2235.830 ;
        RECT 2712.260 2235.170 2712.520 2235.490 ;
        RECT 2712.320 2221.890 2712.460 2235.170 ;
        RECT 2710.880 2221.570 2711.140 2221.890 ;
        RECT 2712.260 2221.570 2712.520 2221.890 ;
        RECT 2710.940 2173.805 2711.080 2221.570 ;
        RECT 2710.870 2173.435 2711.150 2173.805 ;
        RECT 2711.790 2173.435 2712.070 2173.805 ;
        RECT 2711.860 2139.270 2712.000 2173.435 ;
        RECT 2711.800 2138.950 2712.060 2139.270 ;
        RECT 2712.260 2138.610 2712.520 2138.930 ;
        RECT 2712.320 2125.330 2712.460 2138.610 ;
        RECT 2710.880 2125.010 2711.140 2125.330 ;
        RECT 2712.260 2125.010 2712.520 2125.330 ;
        RECT 2710.940 2077.245 2711.080 2125.010 ;
        RECT 2710.870 2076.875 2711.150 2077.245 ;
        RECT 2711.790 2076.875 2712.070 2077.245 ;
        RECT 2711.860 2042.710 2712.000 2076.875 ;
        RECT 2711.800 2042.390 2712.060 2042.710 ;
        RECT 2712.260 2041.710 2712.520 2042.030 ;
        RECT 2712.320 2028.430 2712.460 2041.710 ;
        RECT 2712.260 2028.110 2712.520 2028.430 ;
        RECT 2712.260 1993.770 2712.520 1994.090 ;
        RECT 2712.320 1946.150 2712.460 1993.770 ;
        RECT 2712.260 1945.830 2712.520 1946.150 ;
        RECT 2712.260 1945.150 2712.520 1945.470 ;
        RECT 2712.320 1897.530 2712.460 1945.150 ;
        RECT 2712.260 1897.210 2712.520 1897.530 ;
        RECT 2713.180 1897.210 2713.440 1897.530 ;
        RECT 2713.240 1859.530 2713.380 1897.210 ;
        RECT 2713.240 1859.390 2713.840 1859.530 ;
        RECT 2713.700 1787.710 2713.840 1859.390 ;
        RECT 2713.640 1787.390 2713.900 1787.710 ;
        RECT 2713.640 1766.650 2713.900 1766.970 ;
        RECT 2713.700 1766.370 2713.840 1766.650 ;
        RECT 2713.700 1766.290 2714.300 1766.370 ;
        RECT 2713.700 1766.230 2714.360 1766.290 ;
        RECT 2714.100 1765.970 2714.360 1766.230 ;
        RECT 2714.100 1703.750 2714.360 1704.070 ;
        RECT 2714.160 1657.570 2714.300 1703.750 ;
        RECT 2713.700 1657.430 2714.300 1657.570 ;
        RECT 2713.700 1628.590 2713.840 1657.430 ;
        RECT 2713.180 1628.270 2713.440 1628.590 ;
        RECT 2713.640 1628.270 2713.900 1628.590 ;
        RECT 2713.240 1594.250 2713.380 1628.270 ;
        RECT 2712.720 1593.930 2712.980 1594.250 ;
        RECT 2713.180 1593.930 2713.440 1594.250 ;
        RECT 2712.780 1559.910 2712.920 1593.930 ;
        RECT 2712.720 1559.590 2712.980 1559.910 ;
        RECT 2713.180 1559.590 2713.440 1559.910 ;
        RECT 2713.240 1511.290 2713.380 1559.590 ;
        RECT 2712.260 1510.970 2712.520 1511.290 ;
        RECT 2713.180 1510.970 2713.440 1511.290 ;
        RECT 2712.320 1510.690 2712.460 1510.970 ;
        RECT 2712.320 1510.550 2712.920 1510.690 ;
        RECT 2712.780 1463.090 2712.920 1510.550 ;
        RECT 2712.780 1462.950 2713.380 1463.090 ;
        RECT 2713.240 1449.070 2713.380 1462.950 ;
        RECT 2713.180 1448.750 2713.440 1449.070 ;
        RECT 2712.260 1400.810 2712.520 1401.130 ;
        RECT 2712.320 1366.530 2712.460 1400.810 ;
        RECT 2712.320 1366.390 2713.380 1366.530 ;
        RECT 2713.240 1338.910 2713.380 1366.390 ;
        RECT 2711.800 1338.590 2712.060 1338.910 ;
        RECT 2713.180 1338.590 2713.440 1338.910 ;
        RECT 2711.860 1221.270 2712.000 1338.590 ;
        RECT 2711.800 1220.950 2712.060 1221.270 ;
        RECT 2713.180 1220.950 2713.440 1221.270 ;
        RECT 2713.240 1173.410 2713.380 1220.950 ;
        RECT 2713.240 1173.270 2713.840 1173.410 ;
        RECT 2713.700 1159.390 2713.840 1173.270 ;
        RECT 2712.720 1159.245 2712.980 1159.390 ;
        RECT 2711.790 1158.875 2712.070 1159.245 ;
        RECT 2712.710 1158.875 2712.990 1159.245 ;
        RECT 2713.640 1159.070 2713.900 1159.390 ;
        RECT 2711.860 1111.110 2712.000 1158.875 ;
        RECT 2711.800 1110.790 2712.060 1111.110 ;
        RECT 2713.180 1110.790 2713.440 1111.110 ;
        RECT 2713.240 1076.850 2713.380 1110.790 ;
        RECT 2713.240 1076.710 2713.840 1076.850 ;
        RECT 2713.700 1062.685 2713.840 1076.710 ;
        RECT 2712.710 1062.315 2712.990 1062.685 ;
        RECT 2713.630 1062.315 2713.910 1062.685 ;
        RECT 2712.780 1014.550 2712.920 1062.315 ;
        RECT 2712.720 1014.230 2712.980 1014.550 ;
        RECT 2713.180 1014.230 2713.440 1014.550 ;
        RECT 2713.240 980.210 2713.380 1014.230 ;
        RECT 2713.180 979.890 2713.440 980.210 ;
        RECT 2713.640 979.550 2713.900 979.870 ;
        RECT 2713.700 966.125 2713.840 979.550 ;
        RECT 2712.710 965.755 2712.990 966.125 ;
        RECT 2713.630 965.755 2713.910 966.125 ;
        RECT 2712.780 917.990 2712.920 965.755 ;
        RECT 2712.720 917.670 2712.980 917.990 ;
        RECT 2714.100 917.670 2714.360 917.990 ;
        RECT 2714.160 869.710 2714.300 917.670 ;
        RECT 2713.180 869.390 2713.440 869.710 ;
        RECT 2714.100 869.390 2714.360 869.710 ;
        RECT 2713.240 845.570 2713.380 869.390 ;
        RECT 2711.800 845.250 2712.060 845.570 ;
        RECT 2713.180 845.250 2713.440 845.570 ;
        RECT 2711.860 807.150 2712.000 845.250 ;
        RECT 2711.800 806.830 2712.060 807.150 ;
        RECT 2713.180 806.830 2713.440 807.150 ;
        RECT 2713.240 759.210 2713.380 806.830 ;
        RECT 2711.800 758.890 2712.060 759.210 ;
        RECT 2713.180 758.890 2713.440 759.210 ;
        RECT 2711.860 710.590 2712.000 758.890 ;
        RECT 2711.800 710.270 2712.060 710.590 ;
        RECT 2713.180 710.270 2713.440 710.590 ;
        RECT 2713.240 662.650 2713.380 710.270 ;
        RECT 2711.800 662.330 2712.060 662.650 ;
        RECT 2713.180 662.330 2713.440 662.650 ;
        RECT 2711.860 641.570 2712.000 662.330 ;
        RECT 2711.800 641.250 2712.060 641.570 ;
        RECT 2713.180 641.250 2713.440 641.570 ;
        RECT 2713.240 603.570 2713.380 641.250 ;
        RECT 2713.240 603.430 2713.840 603.570 ;
        RECT 2713.700 579.885 2713.840 603.430 ;
        RECT 2711.800 579.370 2712.060 579.690 ;
        RECT 2712.710 579.515 2712.990 579.885 ;
        RECT 2713.630 579.515 2713.910 579.885 ;
        RECT 2712.720 579.370 2712.980 579.515 ;
        RECT 2711.860 531.605 2712.000 579.370 ;
        RECT 2711.790 531.235 2712.070 531.605 ;
        RECT 2713.170 531.235 2713.450 531.605 ;
        RECT 2713.240 507.270 2713.380 531.235 ;
        RECT 2713.180 506.950 2713.440 507.270 ;
        RECT 2713.640 496.410 2713.900 496.730 ;
        RECT 2713.700 448.530 2713.840 496.410 ;
        RECT 2713.240 448.390 2713.840 448.530 ;
        RECT 2713.240 400.365 2713.380 448.390 ;
        RECT 2713.170 399.995 2713.450 400.365 ;
        RECT 2713.170 386.395 2713.450 386.765 ;
        RECT 2713.240 386.085 2713.380 386.395 ;
        RECT 2713.170 385.715 2713.450 386.085 ;
        RECT 2712.710 338.115 2712.990 338.485 ;
        RECT 2712.780 337.950 2712.920 338.115 ;
        RECT 2712.720 337.630 2712.980 337.950 ;
        RECT 2713.640 337.630 2713.900 337.950 ;
        RECT 2713.700 303.010 2713.840 337.630 ;
        RECT 2713.240 302.870 2713.840 303.010 ;
        RECT 519.850 216.000 520.130 220.000 ;
        RECT 519.960 205.690 520.100 216.000 ;
        RECT 2713.240 210.645 2713.380 302.870 ;
        RECT 607.290 210.275 607.570 210.645 ;
        RECT 2713.170 210.275 2713.450 210.645 ;
        RECT 607.360 205.690 607.500 210.275 ;
        RECT 519.900 205.370 520.160 205.690 ;
        RECT 607.300 205.370 607.560 205.690 ;
      LAYER via2 ;
        RECT 2712.710 2608.000 2712.990 2608.280 ;
        RECT 2713.630 2608.000 2713.910 2608.280 ;
        RECT 2711.790 2511.440 2712.070 2511.720 ;
        RECT 2713.170 2511.440 2713.450 2511.720 ;
        RECT 2711.790 2463.160 2712.070 2463.440 ;
        RECT 2712.710 2463.160 2712.990 2463.440 ;
        RECT 2711.790 2270.040 2712.070 2270.320 ;
        RECT 2713.170 2270.040 2713.450 2270.320 ;
        RECT 2710.870 2173.480 2711.150 2173.760 ;
        RECT 2711.790 2173.480 2712.070 2173.760 ;
        RECT 2710.870 2076.920 2711.150 2077.200 ;
        RECT 2711.790 2076.920 2712.070 2077.200 ;
        RECT 2711.790 1158.920 2712.070 1159.200 ;
        RECT 2712.710 1158.920 2712.990 1159.200 ;
        RECT 2712.710 1062.360 2712.990 1062.640 ;
        RECT 2713.630 1062.360 2713.910 1062.640 ;
        RECT 2712.710 965.800 2712.990 966.080 ;
        RECT 2713.630 965.800 2713.910 966.080 ;
        RECT 2712.710 579.560 2712.990 579.840 ;
        RECT 2713.630 579.560 2713.910 579.840 ;
        RECT 2711.790 531.280 2712.070 531.560 ;
        RECT 2713.170 531.280 2713.450 531.560 ;
        RECT 2713.170 400.040 2713.450 400.320 ;
        RECT 2713.170 386.440 2713.450 386.720 ;
        RECT 2713.170 385.760 2713.450 386.040 ;
        RECT 2712.710 338.160 2712.990 338.440 ;
        RECT 607.290 210.320 607.570 210.600 ;
        RECT 2713.170 210.320 2713.450 210.600 ;
      LAYER met3 ;
        RECT 2712.685 2608.290 2713.015 2608.305 ;
        RECT 2713.605 2608.290 2713.935 2608.305 ;
        RECT 2712.685 2607.990 2713.935 2608.290 ;
        RECT 2712.685 2607.975 2713.015 2607.990 ;
        RECT 2713.605 2607.975 2713.935 2607.990 ;
        RECT 2711.765 2511.730 2712.095 2511.745 ;
        RECT 2713.145 2511.730 2713.475 2511.745 ;
        RECT 2711.765 2511.430 2713.475 2511.730 ;
        RECT 2711.765 2511.415 2712.095 2511.430 ;
        RECT 2713.145 2511.415 2713.475 2511.430 ;
        RECT 2711.765 2463.450 2712.095 2463.465 ;
        RECT 2712.685 2463.450 2713.015 2463.465 ;
        RECT 2711.765 2463.150 2713.015 2463.450 ;
        RECT 2711.765 2463.135 2712.095 2463.150 ;
        RECT 2712.685 2463.135 2713.015 2463.150 ;
        RECT 2711.765 2270.330 2712.095 2270.345 ;
        RECT 2713.145 2270.330 2713.475 2270.345 ;
        RECT 2711.765 2270.030 2713.475 2270.330 ;
        RECT 2711.765 2270.015 2712.095 2270.030 ;
        RECT 2713.145 2270.015 2713.475 2270.030 ;
        RECT 2710.845 2173.770 2711.175 2173.785 ;
        RECT 2711.765 2173.770 2712.095 2173.785 ;
        RECT 2710.845 2173.470 2712.095 2173.770 ;
        RECT 2710.845 2173.455 2711.175 2173.470 ;
        RECT 2711.765 2173.455 2712.095 2173.470 ;
        RECT 2710.845 2077.210 2711.175 2077.225 ;
        RECT 2711.765 2077.210 2712.095 2077.225 ;
        RECT 2710.845 2076.910 2712.095 2077.210 ;
        RECT 2710.845 2076.895 2711.175 2076.910 ;
        RECT 2711.765 2076.895 2712.095 2076.910 ;
        RECT 2711.765 1159.210 2712.095 1159.225 ;
        RECT 2712.685 1159.210 2713.015 1159.225 ;
        RECT 2711.765 1158.910 2713.015 1159.210 ;
        RECT 2711.765 1158.895 2712.095 1158.910 ;
        RECT 2712.685 1158.895 2713.015 1158.910 ;
        RECT 2712.685 1062.650 2713.015 1062.665 ;
        RECT 2713.605 1062.650 2713.935 1062.665 ;
        RECT 2712.685 1062.350 2713.935 1062.650 ;
        RECT 2712.685 1062.335 2713.015 1062.350 ;
        RECT 2713.605 1062.335 2713.935 1062.350 ;
        RECT 2712.685 966.090 2713.015 966.105 ;
        RECT 2713.605 966.090 2713.935 966.105 ;
        RECT 2712.685 965.790 2713.935 966.090 ;
        RECT 2712.685 965.775 2713.015 965.790 ;
        RECT 2713.605 965.775 2713.935 965.790 ;
        RECT 2712.685 579.850 2713.015 579.865 ;
        RECT 2713.605 579.850 2713.935 579.865 ;
        RECT 2712.685 579.550 2713.935 579.850 ;
        RECT 2712.685 579.535 2713.015 579.550 ;
        RECT 2713.605 579.535 2713.935 579.550 ;
        RECT 2711.765 531.570 2712.095 531.585 ;
        RECT 2713.145 531.570 2713.475 531.585 ;
        RECT 2711.765 531.270 2713.475 531.570 ;
        RECT 2711.765 531.255 2712.095 531.270 ;
        RECT 2713.145 531.255 2713.475 531.270 ;
        RECT 2713.145 400.340 2713.475 400.345 ;
        RECT 2713.145 400.330 2713.730 400.340 ;
        RECT 2713.145 400.030 2713.930 400.330 ;
        RECT 2713.145 400.020 2713.730 400.030 ;
        RECT 2713.145 400.015 2713.475 400.020 ;
        RECT 2713.145 386.740 2713.475 386.745 ;
        RECT 2713.145 386.730 2713.730 386.740 ;
        RECT 2713.145 386.430 2713.930 386.730 ;
        RECT 2713.145 386.420 2713.730 386.430 ;
        RECT 2713.145 386.415 2713.475 386.420 ;
        RECT 2712.430 386.050 2712.810 386.060 ;
        RECT 2713.145 386.050 2713.475 386.065 ;
        RECT 2712.430 385.750 2713.475 386.050 ;
        RECT 2712.430 385.740 2712.810 385.750 ;
        RECT 2713.145 385.735 2713.475 385.750 ;
        RECT 2712.685 338.460 2713.015 338.465 ;
        RECT 2712.430 338.450 2713.015 338.460 ;
        RECT 2712.430 338.150 2713.240 338.450 ;
        RECT 2712.430 338.140 2713.015 338.150 ;
        RECT 2712.685 338.135 2713.015 338.140 ;
        RECT 607.265 210.610 607.595 210.625 ;
        RECT 2713.145 210.610 2713.475 210.625 ;
        RECT 607.265 210.310 2713.475 210.610 ;
        RECT 607.265 210.295 607.595 210.310 ;
        RECT 2713.145 210.295 2713.475 210.310 ;
      LAYER via3 ;
        RECT 2713.380 400.020 2713.700 400.340 ;
        RECT 2713.380 386.420 2713.700 386.740 ;
        RECT 2712.460 385.740 2712.780 386.060 ;
        RECT 2712.460 338.140 2712.780 338.460 ;
      LAYER met4 ;
        RECT 2713.375 400.015 2713.705 400.345 ;
        RECT 2713.390 386.745 2713.690 400.015 ;
        RECT 2713.375 386.415 2713.705 386.745 ;
        RECT 2712.455 385.735 2712.785 386.065 ;
        RECT 2712.470 338.465 2712.770 385.735 ;
        RECT 2712.455 338.135 2712.785 338.465 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1997.390 3501.560 1997.710 3501.620 ;
        RECT 2392.530 3501.560 2392.850 3501.620 ;
        RECT 1997.390 3501.420 2392.850 3501.560 ;
        RECT 1997.390 3501.360 1997.710 3501.420 ;
        RECT 2392.530 3501.360 2392.850 3501.420 ;
      LAYER via ;
        RECT 1997.420 3501.360 1997.680 3501.620 ;
        RECT 2392.560 3501.360 2392.820 3501.620 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3501.650 2392.760 3517.600 ;
        RECT 1997.420 3501.330 1997.680 3501.650 ;
        RECT 2392.560 3501.330 2392.820 3501.650 ;
        RECT 1029.530 216.000 1029.810 220.000 ;
        RECT 1029.640 212.685 1029.780 216.000 ;
        RECT 1997.480 212.685 1997.620 3501.330 ;
        RECT 1029.570 212.315 1029.850 212.685 ;
        RECT 1997.410 212.315 1997.690 212.685 ;
      LAYER via2 ;
        RECT 1029.570 212.360 1029.850 212.640 ;
        RECT 1997.410 212.360 1997.690 212.640 ;
      LAYER met3 ;
        RECT 1029.545 212.650 1029.875 212.665 ;
        RECT 1997.385 212.650 1997.715 212.665 ;
        RECT 1029.545 212.350 1997.715 212.650 ;
        RECT 1029.545 212.335 1029.875 212.350 ;
        RECT 1997.385 212.335 1997.715 212.350 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1452.290 3501.900 1452.610 3501.960 ;
        RECT 2068.230 3501.900 2068.550 3501.960 ;
        RECT 1452.290 3501.760 2068.550 3501.900 ;
        RECT 1452.290 3501.700 1452.610 3501.760 ;
        RECT 2068.230 3501.700 2068.550 3501.760 ;
        RECT 1419.170 469.100 1419.490 469.160 ;
        RECT 1452.290 469.100 1452.610 469.160 ;
        RECT 1419.170 468.960 1452.610 469.100 ;
        RECT 1419.170 468.900 1419.490 468.960 ;
        RECT 1452.290 468.900 1452.610 468.960 ;
      LAYER via ;
        RECT 1452.320 3501.700 1452.580 3501.960 ;
        RECT 2068.260 3501.700 2068.520 3501.960 ;
        RECT 1419.200 468.900 1419.460 469.160 ;
        RECT 1452.320 468.900 1452.580 469.160 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3501.990 2068.460 3517.600 ;
        RECT 1452.320 3501.670 1452.580 3501.990 ;
        RECT 2068.260 3501.670 2068.520 3501.990 ;
        RECT 1452.380 469.190 1452.520 3501.670 ;
        RECT 1419.200 468.870 1419.460 469.190 ;
        RECT 1452.320 468.870 1452.580 469.190 ;
        RECT 1419.260 468.365 1419.400 468.870 ;
        RECT 1419.190 467.995 1419.470 468.365 ;
      LAYER via2 ;
        RECT 1419.190 468.040 1419.470 468.320 ;
      LAYER met3 ;
        RECT 1419.165 468.330 1419.495 468.345 ;
        RECT 1408.060 468.240 1419.495 468.330 ;
        RECT 1404.305 468.030 1419.495 468.240 ;
        RECT 1404.305 467.640 1408.305 468.030 ;
        RECT 1419.165 468.015 1419.495 468.030 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 717.210 3502.240 717.530 3502.300 ;
        RECT 1743.930 3502.240 1744.250 3502.300 ;
        RECT 717.210 3502.100 1744.250 3502.240 ;
        RECT 717.210 3502.040 717.530 3502.100 ;
        RECT 1743.930 3502.040 1744.250 3502.100 ;
      LAYER via ;
        RECT 717.240 3502.040 717.500 3502.300 ;
        RECT 1743.960 3502.040 1744.220 3502.300 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3502.330 1744.160 3517.600 ;
        RECT 717.240 3502.010 717.500 3502.330 ;
        RECT 1743.960 3502.010 1744.220 3502.330 ;
        RECT 717.300 1325.050 717.440 3502.010 ;
        RECT 715.990 1325.025 717.440 1325.050 ;
        RECT 715.810 1324.910 717.440 1325.025 ;
        RECT 715.810 1321.025 716.090 1324.910 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1414.570 3464.160 1414.890 3464.220 ;
        RECT 1419.170 3464.160 1419.490 3464.220 ;
        RECT 1414.570 3464.020 1419.490 3464.160 ;
        RECT 1414.570 3463.960 1414.890 3464.020 ;
        RECT 1419.170 3463.960 1419.490 3464.020 ;
      LAYER via ;
        RECT 1414.600 3463.960 1414.860 3464.220 ;
        RECT 1419.200 3463.960 1419.460 3464.220 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3464.250 1419.400 3517.600 ;
        RECT 1414.600 3463.930 1414.860 3464.250 ;
        RECT 1419.200 3463.930 1419.460 3464.250 ;
        RECT 1414.660 1187.010 1414.800 3463.930 ;
        RECT 1414.200 1186.870 1414.800 1187.010 ;
        RECT 1414.200 262.325 1414.340 1186.870 ;
        RECT 1414.130 261.955 1414.410 262.325 ;
        RECT 480.290 216.000 480.570 220.000 ;
        RECT 480.400 204.525 480.540 216.000 ;
        RECT 480.330 204.155 480.610 204.525 ;
      LAYER via2 ;
        RECT 1414.130 262.000 1414.410 262.280 ;
        RECT 480.330 204.200 480.610 204.480 ;
      LAYER met3 ;
        RECT 1409.710 262.290 1410.090 262.300 ;
        RECT 1414.105 262.290 1414.435 262.305 ;
        RECT 1409.710 261.990 1414.435 262.290 ;
        RECT 1409.710 261.980 1410.090 261.990 ;
        RECT 1414.105 261.975 1414.435 261.990 ;
        RECT 480.305 204.490 480.635 204.505 ;
        RECT 1409.710 204.490 1410.090 204.500 ;
        RECT 480.305 204.190 1410.090 204.490 ;
        RECT 480.305 204.175 480.635 204.190 ;
        RECT 1409.710 204.180 1410.090 204.190 ;
      LAYER via3 ;
        RECT 1409.740 261.980 1410.060 262.300 ;
        RECT 1409.740 204.180 1410.060 204.500 ;
      LAYER met4 ;
        RECT 1409.735 261.975 1410.065 262.305 ;
        RECT 1409.750 204.505 1410.050 261.975 ;
        RECT 1409.735 204.175 1410.065 204.505 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1101.310 1342.900 1101.630 1342.960 ;
        RECT 1473.450 1342.900 1473.770 1342.960 ;
        RECT 1101.310 1342.760 1473.770 1342.900 ;
        RECT 1101.310 1342.700 1101.630 1342.760 ;
        RECT 1473.450 1342.700 1473.770 1342.760 ;
        RECT 1473.450 386.140 1473.770 386.200 ;
        RECT 2898.070 386.140 2898.390 386.200 ;
        RECT 1473.450 386.000 2898.390 386.140 ;
        RECT 1473.450 385.940 1473.770 386.000 ;
        RECT 2898.070 385.940 2898.390 386.000 ;
      LAYER via ;
        RECT 1101.340 1342.700 1101.600 1342.960 ;
        RECT 1473.480 1342.700 1473.740 1342.960 ;
        RECT 1473.480 385.940 1473.740 386.200 ;
        RECT 2898.100 385.940 2898.360 386.200 ;
      LAYER met2 ;
        RECT 1101.340 1342.670 1101.600 1342.990 ;
        RECT 1473.480 1342.670 1473.740 1342.990 ;
        RECT 1101.400 1325.025 1101.540 1342.670 ;
        RECT 1101.290 1321.025 1101.570 1325.025 ;
        RECT 1473.540 386.230 1473.680 1342.670 ;
        RECT 1473.480 385.910 1473.740 386.230 ;
        RECT 2898.100 385.910 2898.360 386.230 ;
        RECT 2898.160 381.325 2898.300 385.910 ;
        RECT 2898.090 380.955 2898.370 381.325 ;
      LAYER via2 ;
        RECT 2898.090 381.000 2898.370 381.280 ;
      LAYER met3 ;
        RECT 2898.065 381.290 2898.395 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2898.065 380.990 2924.800 381.290 ;
        RECT 2898.065 380.975 2898.395 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3501.845 1095.100 3517.600 ;
        RECT 1094.890 3501.475 1095.170 3501.845 ;
        RECT 500.530 216.000 500.810 220.000 ;
        RECT 500.640 206.565 500.780 216.000 ;
        RECT 500.570 206.195 500.850 206.565 ;
      LAYER via2 ;
        RECT 1094.890 3501.520 1095.170 3501.800 ;
        RECT 500.570 206.240 500.850 206.520 ;
      LAYER met3 ;
        RECT 281.790 3501.810 282.170 3501.820 ;
        RECT 1094.865 3501.810 1095.195 3501.825 ;
        RECT 281.790 3501.510 1095.195 3501.810 ;
        RECT 281.790 3501.500 282.170 3501.510 ;
        RECT 1094.865 3501.495 1095.195 3501.510 ;
        RECT 281.790 206.530 282.170 206.540 ;
        RECT 500.545 206.530 500.875 206.545 ;
        RECT 281.790 206.230 500.875 206.530 ;
        RECT 281.790 206.220 282.170 206.230 ;
        RECT 500.545 206.215 500.875 206.230 ;
      LAYER via3 ;
        RECT 281.820 3501.500 282.140 3501.820 ;
        RECT 281.820 206.220 282.140 206.540 ;
      LAYER met4 ;
        RECT 281.815 3501.495 282.145 3501.825 ;
        RECT 281.830 206.545 282.130 3501.495 ;
        RECT 281.815 206.215 282.145 206.545 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.510 3503.600 558.830 3503.660 ;
        RECT 770.570 3503.600 770.890 3503.660 ;
        RECT 558.510 3503.460 770.890 3503.600 ;
        RECT 558.510 3503.400 558.830 3503.460 ;
        RECT 770.570 3503.400 770.890 3503.460 ;
        RECT 552.070 1338.480 552.390 1338.540 ;
        RECT 558.510 1338.480 558.830 1338.540 ;
        RECT 552.070 1338.340 558.830 1338.480 ;
        RECT 552.070 1338.280 552.390 1338.340 ;
        RECT 558.510 1338.280 558.830 1338.340 ;
      LAYER via ;
        RECT 558.540 3503.400 558.800 3503.660 ;
        RECT 770.600 3503.400 770.860 3503.660 ;
        RECT 552.100 1338.280 552.360 1338.540 ;
        RECT 558.540 1338.280 558.800 1338.540 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3503.690 770.800 3517.600 ;
        RECT 558.540 3503.370 558.800 3503.690 ;
        RECT 770.600 3503.370 770.860 3503.690 ;
        RECT 558.600 1338.570 558.740 3503.370 ;
        RECT 552.100 1338.250 552.360 1338.570 ;
        RECT 558.540 1338.250 558.800 1338.570 ;
        RECT 552.160 1325.025 552.300 1338.250 ;
        RECT 552.050 1321.025 552.330 1325.025 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 1390.160 448.430 1390.220 ;
        RECT 1416.870 1390.160 1417.190 1390.220 ;
        RECT 448.110 1390.020 1417.190 1390.160 ;
        RECT 448.110 1389.960 448.430 1390.020 ;
        RECT 1416.870 1389.960 1417.190 1390.020 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 1389.960 448.400 1390.220 ;
        RECT 1416.900 1389.960 1417.160 1390.220 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 1390.250 448.340 3498.270 ;
        RECT 448.140 1389.930 448.400 1390.250 ;
        RECT 1416.900 1389.930 1417.160 1390.250 ;
        RECT 1416.960 806.210 1417.100 1389.930 ;
        RECT 1416.500 806.070 1417.100 806.210 ;
        RECT 1416.500 782.525 1416.640 806.070 ;
        RECT 1416.430 782.155 1416.710 782.525 ;
      LAYER via2 ;
        RECT 1416.430 782.200 1416.710 782.480 ;
      LAYER met3 ;
        RECT 1416.405 782.490 1416.735 782.505 ;
        RECT 1408.060 782.400 1416.735 782.490 ;
        RECT 1404.305 782.190 1416.735 782.400 ;
        RECT 1404.305 781.800 1408.305 782.190 ;
        RECT 1416.405 782.175 1416.735 782.190 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.900 121.830 3501.960 ;
        RECT 1269.670 3501.900 1269.990 3501.960 ;
        RECT 121.510 3501.760 1269.990 3501.900 ;
        RECT 121.510 3501.700 121.830 3501.760 ;
        RECT 1269.670 3501.700 1269.990 3501.760 ;
      LAYER via ;
        RECT 121.540 3501.700 121.800 3501.960 ;
        RECT 1269.700 3501.700 1269.960 3501.960 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.990 121.740 3517.600 ;
        RECT 121.540 3501.670 121.800 3501.990 ;
        RECT 1269.700 3501.670 1269.960 3501.990 ;
        RECT 1269.760 1325.025 1269.900 3501.670 ;
        RECT 1269.650 1321.025 1269.930 1325.025 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 258.590 3339.720 258.910 3339.780 ;
        RECT 17.090 3339.580 258.910 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 258.590 3339.520 258.910 3339.580 ;
        RECT 258.590 209.680 258.910 209.740 ;
        RECT 1291.750 209.680 1292.070 209.740 ;
        RECT 258.590 209.540 1292.070 209.680 ;
        RECT 258.590 209.480 258.910 209.540 ;
        RECT 1291.750 209.480 1292.070 209.540 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 258.620 3339.520 258.880 3339.780 ;
        RECT 258.620 209.480 258.880 209.740 ;
        RECT 1291.780 209.480 1292.040 209.740 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 258.620 3339.490 258.880 3339.810 ;
        RECT 258.680 209.770 258.820 3339.490 ;
        RECT 1291.730 216.000 1292.010 220.000 ;
        RECT 1291.840 209.770 1291.980 216.000 ;
        RECT 258.620 209.450 258.880 209.770 ;
        RECT 1291.780 209.450 1292.040 209.770 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 72.750 3050.040 73.070 3050.100 ;
        RECT 17.090 3049.900 73.070 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 72.750 3049.840 73.070 3049.900 ;
        RECT 72.750 1083.140 73.070 1083.200 ;
        RECT 296.770 1083.140 297.090 1083.200 ;
        RECT 72.750 1083.000 297.090 1083.140 ;
        RECT 72.750 1082.940 73.070 1083.000 ;
        RECT 296.770 1082.940 297.090 1083.000 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 72.780 3049.840 73.040 3050.100 ;
        RECT 72.780 1082.940 73.040 1083.200 ;
        RECT 296.800 1082.940 297.060 1083.200 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 72.780 3049.810 73.040 3050.130 ;
        RECT 72.840 1083.230 72.980 3049.810 ;
        RECT 72.780 1082.910 73.040 1083.230 ;
        RECT 296.800 1083.085 297.060 1083.230 ;
        RECT 296.790 1082.715 297.070 1083.085 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
        RECT 296.790 1082.760 297.070 1083.040 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
        RECT 296.765 1083.050 297.095 1083.065 ;
        RECT 296.765 1082.960 310.500 1083.050 ;
        RECT 296.765 1082.750 314.000 1082.960 ;
        RECT 296.765 1082.735 297.095 1082.750 ;
        RECT 310.000 1082.360 314.000 1082.750 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 2760.360 20.630 2760.420 ;
        RECT 79.190 2760.360 79.510 2760.420 ;
        RECT 20.310 2760.220 79.510 2760.360 ;
        RECT 20.310 2760.160 20.630 2760.220 ;
        RECT 79.190 2760.160 79.510 2760.220 ;
        RECT 79.190 841.740 79.510 841.800 ;
        RECT 296.770 841.740 297.090 841.800 ;
        RECT 79.190 841.600 297.090 841.740 ;
        RECT 79.190 841.540 79.510 841.600 ;
        RECT 296.770 841.540 297.090 841.600 ;
      LAYER via ;
        RECT 20.340 2760.160 20.600 2760.420 ;
        RECT 79.220 2760.160 79.480 2760.420 ;
        RECT 79.220 841.540 79.480 841.800 ;
        RECT 296.800 841.540 297.060 841.800 ;
      LAYER met2 ;
        RECT 20.330 2765.035 20.610 2765.405 ;
        RECT 20.400 2760.450 20.540 2765.035 ;
        RECT 20.340 2760.130 20.600 2760.450 ;
        RECT 79.220 2760.130 79.480 2760.450 ;
        RECT 79.280 841.830 79.420 2760.130 ;
        RECT 79.220 841.510 79.480 841.830 ;
        RECT 296.800 841.510 297.060 841.830 ;
        RECT 296.860 841.005 297.000 841.510 ;
        RECT 296.790 840.635 297.070 841.005 ;
      LAYER via2 ;
        RECT 20.330 2765.080 20.610 2765.360 ;
        RECT 296.790 840.680 297.070 840.960 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 20.305 2765.370 20.635 2765.385 ;
        RECT -4.800 2765.070 20.635 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 20.305 2765.055 20.635 2765.070 ;
        RECT 296.765 840.970 297.095 840.985 ;
        RECT 296.765 840.880 310.500 840.970 ;
        RECT 296.765 840.670 314.000 840.880 ;
        RECT 296.765 840.655 297.095 840.670 ;
        RECT 310.000 840.280 314.000 840.670 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 2477.480 20.630 2477.540 ;
        RECT 1028.170 2477.480 1028.490 2477.540 ;
        RECT 20.310 2477.340 1028.490 2477.480 ;
        RECT 20.310 2477.280 20.630 2477.340 ;
        RECT 1028.170 2477.280 1028.490 2477.340 ;
      LAYER via ;
        RECT 20.340 2477.280 20.600 2477.540 ;
        RECT 1028.200 2477.280 1028.460 2477.540 ;
      LAYER met2 ;
        RECT 20.330 2477.395 20.610 2477.765 ;
        RECT 20.340 2477.250 20.600 2477.395 ;
        RECT 1028.200 2477.250 1028.460 2477.570 ;
        RECT 1028.260 1337.290 1028.400 2477.250 ;
        RECT 1028.260 1337.150 1030.700 1337.290 ;
        RECT 1030.560 1325.050 1030.700 1337.150 ;
        RECT 1030.560 1325.025 1032.470 1325.050 ;
        RECT 1030.560 1324.910 1032.570 1325.025 ;
        RECT 1032.290 1321.025 1032.570 1324.910 ;
      LAYER via2 ;
        RECT 20.330 2477.440 20.610 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 20.305 2477.730 20.635 2477.745 ;
        RECT -4.800 2477.430 20.635 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 20.305 2477.415 20.635 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.930 2187.460 19.250 2187.520 ;
        RECT 72.290 2187.460 72.610 2187.520 ;
        RECT 18.930 2187.320 72.610 2187.460 ;
        RECT 18.930 2187.260 19.250 2187.320 ;
        RECT 72.290 2187.260 72.610 2187.320 ;
        RECT 72.290 199.820 72.610 199.880 ;
        RECT 1321.190 199.820 1321.510 199.880 ;
        RECT 72.290 199.680 1321.510 199.820 ;
        RECT 72.290 199.620 72.610 199.680 ;
        RECT 1321.190 199.620 1321.510 199.680 ;
      LAYER via ;
        RECT 18.960 2187.260 19.220 2187.520 ;
        RECT 72.320 2187.260 72.580 2187.520 ;
        RECT 72.320 199.620 72.580 199.880 ;
        RECT 1321.220 199.620 1321.480 199.880 ;
      LAYER met2 ;
        RECT 18.950 2189.755 19.230 2190.125 ;
        RECT 19.020 2187.550 19.160 2189.755 ;
        RECT 18.960 2187.230 19.220 2187.550 ;
        RECT 72.320 2187.230 72.580 2187.550 ;
        RECT 72.380 199.910 72.520 2187.230 ;
        RECT 1321.170 216.000 1321.450 220.000 ;
        RECT 1321.280 199.910 1321.420 216.000 ;
        RECT 72.320 199.590 72.580 199.910 ;
        RECT 1321.220 199.590 1321.480 199.910 ;
      LAYER via2 ;
        RECT 18.950 2189.800 19.230 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 18.925 2190.090 19.255 2190.105 ;
        RECT -4.800 2189.790 19.255 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 18.925 2189.775 19.255 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 19.850 1897.780 20.170 1897.840 ;
        RECT 120.590 1897.780 120.910 1897.840 ;
        RECT 19.850 1897.640 120.910 1897.780 ;
        RECT 19.850 1897.580 20.170 1897.640 ;
        RECT 120.590 1897.580 120.910 1897.640 ;
        RECT 120.590 1000.520 120.910 1000.580 ;
        RECT 296.770 1000.520 297.090 1000.580 ;
        RECT 120.590 1000.380 297.090 1000.520 ;
        RECT 120.590 1000.320 120.910 1000.380 ;
        RECT 296.770 1000.320 297.090 1000.380 ;
      LAYER via ;
        RECT 19.880 1897.580 20.140 1897.840 ;
        RECT 120.620 1897.580 120.880 1897.840 ;
        RECT 120.620 1000.320 120.880 1000.580 ;
        RECT 296.800 1000.320 297.060 1000.580 ;
      LAYER met2 ;
        RECT 19.870 1902.795 20.150 1903.165 ;
        RECT 19.940 1897.870 20.080 1902.795 ;
        RECT 19.880 1897.550 20.140 1897.870 ;
        RECT 120.620 1897.550 120.880 1897.870 ;
        RECT 120.680 1000.610 120.820 1897.550 ;
        RECT 120.620 1000.290 120.880 1000.610 ;
        RECT 296.800 1000.290 297.060 1000.610 ;
        RECT 296.860 994.685 297.000 1000.290 ;
        RECT 296.790 994.315 297.070 994.685 ;
      LAYER via2 ;
        RECT 19.870 1902.840 20.150 1903.120 ;
        RECT 296.790 994.360 297.070 994.640 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 19.845 1903.130 20.175 1903.145 ;
        RECT -4.800 1902.830 20.175 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 19.845 1902.815 20.175 1902.830 ;
        RECT 296.765 994.650 297.095 994.665 ;
        RECT 296.765 994.560 310.500 994.650 ;
        RECT 296.765 994.350 314.000 994.560 ;
        RECT 296.765 994.335 297.095 994.350 ;
        RECT 310.000 993.960 314.000 994.350 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1420.090 766.260 1420.410 766.320 ;
        RECT 1611.450 766.260 1611.770 766.320 ;
        RECT 1420.090 766.120 1611.770 766.260 ;
        RECT 1420.090 766.060 1420.410 766.120 ;
        RECT 1611.450 766.060 1611.770 766.120 ;
        RECT 1611.450 620.740 1611.770 620.800 ;
        RECT 2899.450 620.740 2899.770 620.800 ;
        RECT 1611.450 620.600 2899.770 620.740 ;
        RECT 1611.450 620.540 1611.770 620.600 ;
        RECT 2899.450 620.540 2899.770 620.600 ;
      LAYER via ;
        RECT 1420.120 766.060 1420.380 766.320 ;
        RECT 1611.480 766.060 1611.740 766.320 ;
        RECT 1611.480 620.540 1611.740 620.800 ;
        RECT 2899.480 620.540 2899.740 620.800 ;
      LAYER met2 ;
        RECT 1420.110 768.555 1420.390 768.925 ;
        RECT 1420.180 766.350 1420.320 768.555 ;
        RECT 1420.120 766.030 1420.380 766.350 ;
        RECT 1611.480 766.030 1611.740 766.350 ;
        RECT 1611.540 620.830 1611.680 766.030 ;
        RECT 1611.480 620.510 1611.740 620.830 ;
        RECT 2899.480 620.510 2899.740 620.830 ;
        RECT 2899.540 615.925 2899.680 620.510 ;
        RECT 2899.470 615.555 2899.750 615.925 ;
      LAYER via2 ;
        RECT 1420.110 768.600 1420.390 768.880 ;
        RECT 2899.470 615.600 2899.750 615.880 ;
      LAYER met3 ;
        RECT 1420.085 768.890 1420.415 768.905 ;
        RECT 1408.060 768.800 1420.415 768.890 ;
        RECT 1404.305 768.590 1420.415 768.800 ;
        RECT 1404.305 768.200 1408.305 768.590 ;
        RECT 1420.085 768.575 1420.415 768.590 ;
        RECT 2899.445 615.890 2899.775 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2899.445 615.590 2924.800 615.890 ;
        RECT 2899.445 615.575 2899.775 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 1117.820 18.330 1117.880 ;
        RECT 296.770 1117.820 297.090 1117.880 ;
        RECT 18.010 1117.680 297.090 1117.820 ;
        RECT 18.010 1117.620 18.330 1117.680 ;
        RECT 296.770 1117.620 297.090 1117.680 ;
      LAYER via ;
        RECT 18.040 1117.620 18.300 1117.880 ;
        RECT 296.800 1117.620 297.060 1117.880 ;
      LAYER met2 ;
        RECT 18.030 1615.155 18.310 1615.525 ;
        RECT 18.100 1117.910 18.240 1615.155 ;
        RECT 18.040 1117.590 18.300 1117.910 ;
        RECT 296.800 1117.590 297.060 1117.910 ;
        RECT 296.860 1111.645 297.000 1117.590 ;
        RECT 296.790 1111.275 297.070 1111.645 ;
      LAYER via2 ;
        RECT 18.030 1615.200 18.310 1615.480 ;
        RECT 296.790 1111.320 297.070 1111.600 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 18.005 1615.490 18.335 1615.505 ;
        RECT -4.800 1615.190 18.335 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 18.005 1615.175 18.335 1615.190 ;
        RECT 296.765 1111.610 297.095 1111.625 ;
        RECT 296.765 1111.520 310.500 1111.610 ;
        RECT 296.765 1111.310 314.000 1111.520 ;
        RECT 296.765 1111.295 297.095 1111.310 ;
        RECT 310.000 1110.920 314.000 1111.310 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.470 945.100 18.790 945.160 ;
        RECT 296.770 945.100 297.090 945.160 ;
        RECT 18.470 944.960 297.090 945.100 ;
        RECT 18.470 944.900 18.790 944.960 ;
        RECT 296.770 944.900 297.090 944.960 ;
      LAYER via ;
        RECT 18.500 944.900 18.760 945.160 ;
        RECT 296.800 944.900 297.060 945.160 ;
      LAYER met2 ;
        RECT 18.490 1400.275 18.770 1400.645 ;
        RECT 18.560 945.190 18.700 1400.275 ;
        RECT 18.500 944.870 18.760 945.190 ;
        RECT 296.800 944.870 297.060 945.190 ;
        RECT 296.860 944.365 297.000 944.870 ;
        RECT 296.790 943.995 297.070 944.365 ;
      LAYER via2 ;
        RECT 18.490 1400.320 18.770 1400.600 ;
        RECT 296.790 944.040 297.070 944.320 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 18.465 1400.610 18.795 1400.625 ;
        RECT -4.800 1400.310 18.795 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 18.465 1400.295 18.795 1400.310 ;
        RECT 296.765 944.330 297.095 944.345 ;
        RECT 296.765 944.240 310.500 944.330 ;
        RECT 296.765 944.030 314.000 944.240 ;
        RECT 296.765 944.015 297.095 944.030 ;
        RECT 310.000 943.640 314.000 944.030 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 86.090 1333.040 86.410 1333.100 ;
        RECT 587.030 1333.040 587.350 1333.100 ;
        RECT 86.090 1332.900 587.350 1333.040 ;
        RECT 86.090 1332.840 86.410 1332.900 ;
        RECT 587.030 1332.840 587.350 1332.900 ;
        RECT 20.310 1186.840 20.630 1186.900 ;
        RECT 86.090 1186.840 86.410 1186.900 ;
        RECT 20.310 1186.700 86.410 1186.840 ;
        RECT 20.310 1186.640 20.630 1186.700 ;
        RECT 86.090 1186.640 86.410 1186.700 ;
      LAYER via ;
        RECT 86.120 1332.840 86.380 1333.100 ;
        RECT 587.060 1332.840 587.320 1333.100 ;
        RECT 20.340 1186.640 20.600 1186.900 ;
        RECT 86.120 1186.640 86.380 1186.900 ;
      LAYER met2 ;
        RECT 86.120 1332.810 86.380 1333.130 ;
        RECT 587.060 1332.810 587.320 1333.130 ;
        RECT 86.180 1186.930 86.320 1332.810 ;
        RECT 587.120 1325.025 587.260 1332.810 ;
        RECT 587.010 1321.025 587.290 1325.025 ;
        RECT 20.340 1186.610 20.600 1186.930 ;
        RECT 86.120 1186.610 86.380 1186.930 ;
        RECT 20.400 1185.085 20.540 1186.610 ;
        RECT 20.330 1184.715 20.610 1185.085 ;
      LAYER via2 ;
        RECT 20.330 1184.760 20.610 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 20.305 1185.050 20.635 1185.065 ;
        RECT -4.800 1184.750 20.635 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 20.305 1184.735 20.635 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 138.070 972.640 138.390 972.700 ;
        RECT 185.910 972.640 186.230 972.700 ;
        RECT 138.070 972.500 186.230 972.640 ;
        RECT 138.070 972.440 138.390 972.500 ;
        RECT 185.910 972.440 186.230 972.500 ;
      LAYER via ;
        RECT 138.100 972.440 138.360 972.700 ;
        RECT 185.940 972.440 186.200 972.700 ;
      LAYER met2 ;
        RECT 1419.190 1173.835 1419.470 1174.205 ;
        RECT 1419.260 1160.605 1419.400 1173.835 ;
        RECT 1419.190 1160.235 1419.470 1160.605 ;
        RECT 24.470 972.555 24.750 972.925 ;
        RECT 61.730 972.555 62.010 972.925 ;
        RECT 110.950 972.555 111.230 972.925 ;
        RECT 138.090 972.555 138.370 972.925 ;
        RECT 24.540 969.525 24.680 972.555 ;
        RECT 61.800 972.130 61.940 972.555 ;
        RECT 62.650 972.130 62.930 972.245 ;
        RECT 61.800 971.990 62.930 972.130 ;
        RECT 62.650 971.875 62.930 971.990 ;
        RECT 110.030 972.130 110.310 972.245 ;
        RECT 111.020 972.130 111.160 972.555 ;
        RECT 138.100 972.410 138.360 972.555 ;
        RECT 185.940 972.410 186.200 972.730 ;
        RECT 110.030 971.990 111.160 972.130 ;
        RECT 110.030 971.875 110.310 971.990 ;
        RECT 186.000 971.565 186.140 972.410 ;
        RECT 185.930 971.195 186.210 971.565 ;
        RECT 24.470 969.155 24.750 969.525 ;
      LAYER via2 ;
        RECT 1419.190 1173.880 1419.470 1174.160 ;
        RECT 1419.190 1160.280 1419.470 1160.560 ;
        RECT 24.470 972.600 24.750 972.880 ;
        RECT 61.730 972.600 62.010 972.880 ;
        RECT 110.950 972.600 111.230 972.880 ;
        RECT 138.090 972.600 138.370 972.880 ;
        RECT 62.650 971.920 62.930 972.200 ;
        RECT 110.030 971.920 110.310 972.200 ;
        RECT 185.930 971.240 186.210 971.520 ;
        RECT 24.470 969.200 24.750 969.480 ;
      LAYER met3 ;
        RECT 1419.165 1174.170 1419.495 1174.185 ;
        RECT 1419.830 1174.170 1420.210 1174.180 ;
        RECT 1419.165 1173.870 1420.210 1174.170 ;
        RECT 1419.165 1173.855 1419.495 1173.870 ;
        RECT 1419.830 1173.860 1420.210 1173.870 ;
        RECT 1419.165 1160.580 1419.495 1160.585 ;
        RECT 1418.910 1160.570 1419.495 1160.580 ;
        RECT 1418.710 1160.270 1419.495 1160.570 ;
        RECT 1418.910 1160.260 1419.495 1160.270 ;
        RECT 1419.165 1160.255 1419.495 1160.260 ;
        RECT 1417.990 1047.010 1418.370 1047.020 ;
        RECT 1407.910 1046.710 1418.370 1047.010 ;
        RECT 1407.910 1046.240 1408.210 1046.710 ;
        RECT 1417.990 1046.700 1418.370 1046.710 ;
        RECT 1404.305 1045.640 1408.305 1046.240 ;
        RECT 24.445 972.890 24.775 972.905 ;
        RECT 61.705 972.890 62.035 972.905 ;
        RECT 24.445 972.590 62.035 972.890 ;
        RECT 24.445 972.575 24.775 972.590 ;
        RECT 61.705 972.575 62.035 972.590 ;
        RECT 110.925 972.890 111.255 972.905 ;
        RECT 138.065 972.890 138.395 972.905 ;
        RECT 110.925 972.590 138.395 972.890 ;
        RECT 110.925 972.575 111.255 972.590 ;
        RECT 138.065 972.575 138.395 972.590 ;
        RECT 275.390 972.590 290.410 972.890 ;
        RECT 62.625 972.210 62.955 972.225 ;
        RECT 110.005 972.210 110.335 972.225 ;
        RECT 275.390 972.210 275.690 972.590 ;
        RECT 62.625 971.910 110.335 972.210 ;
        RECT 62.625 971.895 62.955 971.910 ;
        RECT 110.005 971.895 110.335 971.910 ;
        RECT 227.550 971.910 275.690 972.210 ;
        RECT 185.905 971.530 186.235 971.545 ;
        RECT 227.550 971.530 227.850 971.910 ;
        RECT 185.905 971.230 227.850 971.530 ;
        RECT 290.110 971.530 290.410 972.590 ;
        RECT 304.790 971.530 305.170 971.540 ;
        RECT 290.110 971.230 305.170 971.530 ;
        RECT 185.905 971.215 186.235 971.230 ;
        RECT 304.790 971.220 305.170 971.230 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 24.445 969.490 24.775 969.505 ;
        RECT -4.800 969.190 24.775 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 24.445 969.175 24.775 969.190 ;
      LAYER via3 ;
        RECT 1419.860 1173.860 1420.180 1174.180 ;
        RECT 1418.940 1160.260 1419.260 1160.580 ;
        RECT 1418.020 1046.700 1418.340 1047.020 ;
        RECT 304.820 971.220 305.140 971.540 ;
      LAYER met4 ;
        RECT 1419.430 1252.310 1420.610 1253.490 ;
        RECT 304.390 1245.510 305.570 1246.690 ;
        RECT 304.830 971.545 305.130 1245.510 ;
        RECT 1419.870 1174.185 1420.170 1252.310 ;
        RECT 1419.855 1173.855 1420.185 1174.185 ;
        RECT 1418.935 1160.255 1419.265 1160.585 ;
        RECT 1418.950 1100.050 1419.250 1160.255 ;
        RECT 1418.030 1099.750 1419.250 1100.050 ;
        RECT 1418.030 1047.025 1418.330 1099.750 ;
        RECT 1418.015 1046.695 1418.345 1047.025 ;
        RECT 304.815 971.215 305.145 971.545 ;
      LAYER met5 ;
        RECT 385.140 1255.500 421.700 1257.100 ;
        RECT 337.300 1248.700 373.860 1250.300 ;
        RECT 337.300 1246.900 338.900 1248.700 ;
        RECT 304.180 1245.300 338.900 1246.900 ;
        RECT 372.260 1246.900 373.860 1248.700 ;
        RECT 385.140 1246.900 386.740 1255.500 ;
        RECT 420.100 1250.300 421.700 1255.500 ;
        RECT 499.220 1255.500 504.500 1257.100 ;
        RECT 499.220 1253.700 500.820 1255.500 ;
        RECT 453.220 1252.100 462.180 1253.700 ;
        RECT 453.220 1250.300 454.820 1252.100 ;
        RECT 420.100 1248.700 454.820 1250.300 ;
        RECT 460.580 1250.300 462.180 1252.100 ;
        RECT 467.940 1252.100 500.820 1253.700 ;
        RECT 502.900 1253.700 504.500 1255.500 ;
        RECT 520.380 1255.500 556.020 1257.100 ;
        RECT 520.380 1253.700 521.980 1255.500 ;
        RECT 502.900 1252.100 521.980 1253.700 ;
        RECT 554.420 1253.700 556.020 1255.500 ;
        RECT 752.220 1255.500 795.220 1257.100 ;
        RECT 554.420 1252.100 558.780 1253.700 ;
        RECT 467.940 1250.300 469.540 1252.100 ;
        RECT 460.580 1248.700 469.540 1250.300 ;
        RECT 557.180 1250.300 558.780 1252.100 ;
        RECT 605.020 1252.100 645.260 1253.700 ;
        RECT 605.020 1250.300 606.620 1252.100 ;
        RECT 557.180 1248.700 561.540 1250.300 ;
        RECT 372.260 1245.300 386.740 1246.900 ;
        RECT 559.940 1246.900 561.540 1248.700 ;
        RECT 584.780 1248.700 606.620 1250.300 ;
        RECT 643.660 1250.300 645.260 1252.100 ;
        RECT 701.620 1252.100 740.020 1253.700 ;
        RECT 701.620 1250.300 703.220 1252.100 ;
        RECT 643.660 1248.700 658.140 1250.300 ;
        RECT 584.780 1246.900 586.380 1248.700 ;
        RECT 559.940 1245.300 586.380 1246.900 ;
        RECT 656.540 1246.900 658.140 1248.700 ;
        RECT 681.380 1248.700 703.220 1250.300 ;
        RECT 681.380 1246.900 682.980 1248.700 ;
        RECT 656.540 1245.300 682.980 1246.900 ;
        RECT 738.420 1246.900 740.020 1252.100 ;
        RECT 752.220 1246.900 753.820 1255.500 ;
        RECT 793.620 1253.700 795.220 1255.500 ;
        RECT 848.820 1255.500 891.820 1257.100 ;
        RECT 793.620 1252.100 836.620 1253.700 ;
        RECT 738.420 1245.300 753.820 1246.900 ;
        RECT 835.020 1246.900 836.620 1252.100 ;
        RECT 848.820 1246.900 850.420 1255.500 ;
        RECT 890.220 1253.700 891.820 1255.500 ;
        RECT 1053.060 1255.500 1077.660 1257.100 ;
        RECT 890.220 1252.100 899.180 1253.700 ;
        RECT 897.580 1250.300 899.180 1252.100 ;
        RECT 946.340 1252.100 984.740 1253.700 ;
        RECT 946.340 1250.300 947.940 1252.100 ;
        RECT 897.580 1248.700 947.940 1250.300 ;
        RECT 835.020 1245.300 850.420 1246.900 ;
        RECT 983.140 1246.900 984.740 1252.100 ;
        RECT 1047.540 1250.300 1050.060 1253.700 ;
        RECT 1053.060 1250.300 1054.660 1255.500 ;
        RECT 1047.540 1248.700 1054.660 1250.300 ;
        RECT 1076.060 1250.300 1077.660 1255.500 ;
        RECT 1149.660 1255.500 1174.260 1257.100 ;
        RECT 1111.020 1252.100 1146.660 1253.700 ;
        RECT 1111.020 1250.300 1112.620 1252.100 ;
        RECT 1076.060 1248.700 1096.980 1250.300 ;
        RECT 1047.540 1246.900 1049.140 1248.700 ;
        RECT 983.140 1245.300 1049.140 1246.900 ;
        RECT 1095.380 1246.900 1096.980 1248.700 ;
        RECT 1110.100 1248.700 1112.620 1250.300 ;
        RECT 1145.060 1250.300 1146.660 1252.100 ;
        RECT 1149.660 1250.300 1151.260 1255.500 ;
        RECT 1145.060 1248.700 1151.260 1250.300 ;
        RECT 1172.660 1250.300 1174.260 1255.500 ;
        RECT 1246.260 1255.500 1270.860 1257.100 ;
        RECT 1207.620 1252.100 1243.260 1253.700 ;
        RECT 1207.620 1250.300 1209.220 1252.100 ;
        RECT 1172.660 1248.700 1193.580 1250.300 ;
        RECT 1110.100 1246.900 1111.700 1248.700 ;
        RECT 1095.380 1245.300 1111.700 1246.900 ;
        RECT 1191.980 1246.900 1193.580 1248.700 ;
        RECT 1206.700 1248.700 1209.220 1250.300 ;
        RECT 1241.660 1250.300 1243.260 1252.100 ;
        RECT 1246.260 1250.300 1247.860 1255.500 ;
        RECT 1241.660 1248.700 1247.860 1250.300 ;
        RECT 1269.260 1250.300 1270.860 1255.500 ;
        RECT 1365.860 1252.100 1420.820 1253.700 ;
        RECT 1365.860 1250.300 1367.460 1252.100 ;
        RECT 1269.260 1248.700 1290.180 1250.300 ;
        RECT 1206.700 1246.900 1208.300 1248.700 ;
        RECT 1191.980 1245.300 1208.300 1246.900 ;
        RECT 1288.580 1246.900 1290.180 1248.700 ;
        RECT 1314.340 1248.700 1367.460 1250.300 ;
        RECT 1314.340 1246.900 1315.940 1248.700 ;
        RECT 1288.580 1245.300 1315.940 1246.900 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 205.260 18.330 205.320 ;
        RECT 534.590 205.260 534.910 205.320 ;
        RECT 18.010 205.120 534.910 205.260 ;
        RECT 18.010 205.060 18.330 205.120 ;
        RECT 534.590 205.060 534.910 205.120 ;
      LAYER via ;
        RECT 18.040 205.060 18.300 205.320 ;
        RECT 534.620 205.060 534.880 205.320 ;
      LAYER met2 ;
        RECT 18.030 753.595 18.310 753.965 ;
        RECT 18.100 205.350 18.240 753.595 ;
        RECT 534.570 216.000 534.850 220.000 ;
        RECT 534.680 205.350 534.820 216.000 ;
        RECT 18.040 205.030 18.300 205.350 ;
        RECT 534.620 205.030 534.880 205.350 ;
      LAYER via2 ;
        RECT 18.030 753.640 18.310 753.920 ;
      LAYER met3 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 18.005 753.930 18.335 753.945 ;
        RECT -4.800 753.630 18.335 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 18.005 753.615 18.335 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 538.460 20.630 538.520 ;
        RECT 278.830 538.460 279.150 538.520 ;
        RECT 20.310 538.320 279.150 538.460 ;
        RECT 20.310 538.260 20.630 538.320 ;
        RECT 278.830 538.260 279.150 538.320 ;
        RECT 278.830 213.080 279.150 213.140 ;
        RECT 802.310 213.080 802.630 213.140 ;
        RECT 278.830 212.940 802.630 213.080 ;
        RECT 278.830 212.880 279.150 212.940 ;
        RECT 802.310 212.880 802.630 212.940 ;
      LAYER via ;
        RECT 20.340 538.260 20.600 538.520 ;
        RECT 278.860 538.260 279.120 538.520 ;
        RECT 278.860 212.880 279.120 213.140 ;
        RECT 802.340 212.880 802.600 213.140 ;
      LAYER met2 ;
        RECT 20.340 538.405 20.600 538.550 ;
        RECT 20.330 538.035 20.610 538.405 ;
        RECT 278.860 538.230 279.120 538.550 ;
        RECT 278.920 213.170 279.060 538.230 ;
        RECT 802.290 216.000 802.570 220.000 ;
        RECT 802.400 213.170 802.540 216.000 ;
        RECT 278.860 212.850 279.120 213.170 ;
        RECT 802.340 212.850 802.600 213.170 ;
      LAYER via2 ;
        RECT 20.330 538.080 20.610 538.360 ;
      LAYER met3 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 20.305 538.370 20.635 538.385 ;
        RECT -4.800 538.070 20.635 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 20.305 538.055 20.635 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 820.710 1334.060 821.030 1334.120 ;
        RECT 987.230 1334.060 987.550 1334.120 ;
        RECT 820.710 1333.920 987.550 1334.060 ;
        RECT 820.710 1333.860 821.030 1333.920 ;
        RECT 987.230 1333.860 987.550 1333.920 ;
        RECT 17.550 1328.620 17.870 1328.680 ;
        RECT 820.710 1328.620 821.030 1328.680 ;
        RECT 17.550 1328.480 821.030 1328.620 ;
        RECT 17.550 1328.420 17.870 1328.480 ;
        RECT 820.710 1328.420 821.030 1328.480 ;
      LAYER via ;
        RECT 820.740 1333.860 821.000 1334.120 ;
        RECT 987.260 1333.860 987.520 1334.120 ;
        RECT 17.580 1328.420 17.840 1328.680 ;
        RECT 820.740 1328.420 821.000 1328.680 ;
      LAYER met2 ;
        RECT 820.740 1333.830 821.000 1334.150 ;
        RECT 987.260 1333.830 987.520 1334.150 ;
        RECT 820.800 1328.710 820.940 1333.830 ;
        RECT 17.580 1328.390 17.840 1328.710 ;
        RECT 820.740 1328.390 821.000 1328.710 ;
        RECT 17.640 322.845 17.780 1328.390 ;
        RECT 987.320 1325.025 987.460 1333.830 ;
        RECT 987.210 1321.025 987.490 1325.025 ;
        RECT 17.570 322.475 17.850 322.845 ;
      LAYER via2 ;
        RECT 17.570 322.520 17.850 322.800 ;
      LAYER met3 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 17.545 322.810 17.875 322.825 ;
        RECT -4.800 322.510 17.875 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 17.545 322.495 17.875 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 732.925 144.925 733.095 168.895 ;
      LAYER mcon ;
        RECT 732.925 168.725 733.095 168.895 ;
      LAYER met1 ;
        RECT 732.850 168.880 733.170 168.940 ;
        RECT 732.655 168.740 733.170 168.880 ;
        RECT 732.850 168.680 733.170 168.740 ;
        RECT 732.865 145.080 733.155 145.125 ;
        RECT 733.310 145.080 733.630 145.140 ;
        RECT 732.865 144.940 733.630 145.080 ;
        RECT 732.865 144.895 733.155 144.940 ;
        RECT 733.310 144.880 733.630 144.940 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 733.310 110.400 733.630 110.460 ;
        RECT 15.710 110.260 733.630 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 733.310 110.200 733.630 110.260 ;
      LAYER via ;
        RECT 732.880 168.680 733.140 168.940 ;
        RECT 733.340 144.880 733.600 145.140 ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 733.340 110.200 733.600 110.460 ;
      LAYER met2 ;
        RECT 737.890 216.650 738.170 220.000 ;
        RECT 732.940 216.510 738.170 216.650 ;
        RECT 732.940 168.970 733.080 216.510 ;
        RECT 737.890 216.000 738.170 216.510 ;
        RECT 732.880 168.650 733.140 168.970 ;
        RECT 733.340 144.850 733.600 145.170 ;
        RECT 733.400 110.490 733.540 144.850 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 733.340 110.170 733.600 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1426.530 848.880 1426.850 848.940 ;
        RECT 2900.830 848.880 2901.150 848.940 ;
        RECT 1426.530 848.740 2901.150 848.880 ;
        RECT 1426.530 848.680 1426.850 848.740 ;
        RECT 2900.830 848.680 2901.150 848.740 ;
        RECT 1277.030 210.020 1277.350 210.080 ;
        RECT 1426.530 210.020 1426.850 210.080 ;
        RECT 1277.030 209.880 1426.850 210.020 ;
        RECT 1277.030 209.820 1277.350 209.880 ;
        RECT 1426.530 209.820 1426.850 209.880 ;
      LAYER via ;
        RECT 1426.560 848.680 1426.820 848.940 ;
        RECT 2900.860 848.680 2901.120 848.940 ;
        RECT 1277.060 209.820 1277.320 210.080 ;
        RECT 1426.560 209.820 1426.820 210.080 ;
      LAYER met2 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
        RECT 2900.920 848.970 2901.060 850.155 ;
        RECT 1426.560 848.650 1426.820 848.970 ;
        RECT 2900.860 848.650 2901.120 848.970 ;
        RECT 1277.010 216.000 1277.290 220.000 ;
        RECT 1277.120 210.110 1277.260 216.000 ;
        RECT 1426.620 210.110 1426.760 848.650 ;
        RECT 1277.060 209.790 1277.320 210.110 ;
        RECT 1426.560 209.790 1426.820 210.110 ;
      LAYER via2 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2903.790 1085.090 2904.170 1085.100 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2903.790 1084.790 2924.800 1085.090 ;
        RECT 2903.790 1084.780 2904.170 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
        RECT 2474.150 386.050 2474.530 386.060 ;
        RECT 2503.590 386.050 2503.970 386.060 ;
        RECT 2474.150 385.750 2503.970 386.050 ;
        RECT 2474.150 385.740 2474.530 385.750 ;
        RECT 2503.590 385.740 2503.970 385.750 ;
        RECT 311.230 382.340 311.610 382.660 ;
        RECT 1406.950 382.650 1407.330 382.660 ;
        RECT 1489.750 382.650 1490.130 382.660 ;
        RECT 1406.950 382.350 1490.130 382.650 ;
        RECT 1406.950 382.340 1407.330 382.350 ;
        RECT 1489.750 382.340 1490.130 382.350 ;
        RECT 1883.510 382.650 1883.890 382.660 ;
        RECT 1948.830 382.650 1949.210 382.660 ;
        RECT 1883.510 382.350 1949.210 382.650 ;
        RECT 1883.510 382.340 1883.890 382.350 ;
        RECT 1948.830 382.340 1949.210 382.350 ;
        RECT 311.270 381.200 311.570 382.340 ;
        RECT 310.000 380.600 314.000 381.200 ;
        RECT 1739.070 379.250 1739.450 379.260 ;
        RECT 1785.990 379.250 1786.370 379.260 ;
        RECT 1739.070 378.950 1786.370 379.250 ;
        RECT 1739.070 378.940 1739.450 378.950 ;
        RECT 1785.990 378.940 1786.370 378.950 ;
      LAYER via3 ;
        RECT 2903.820 1084.780 2904.140 1085.100 ;
        RECT 2474.180 385.740 2474.500 386.060 ;
        RECT 2503.620 385.740 2503.940 386.060 ;
        RECT 311.260 382.340 311.580 382.660 ;
        RECT 1406.980 382.340 1407.300 382.660 ;
        RECT 1489.780 382.340 1490.100 382.660 ;
        RECT 1883.540 382.340 1883.860 382.660 ;
        RECT 1948.860 382.340 1949.180 382.660 ;
        RECT 1739.100 378.940 1739.420 379.260 ;
        RECT 1786.020 378.940 1786.340 379.260 ;
      LAYER met4 ;
        RECT 2903.815 1084.775 2904.145 1085.105 ;
        RECT 1489.350 385.310 1490.530 386.490 ;
        RECT 2473.750 385.310 2474.930 386.490 ;
        RECT 2503.615 385.735 2503.945 386.065 ;
        RECT 310.830 381.910 312.010 383.090 ;
        RECT 1406.550 381.910 1407.730 383.090 ;
        RECT 1489.790 382.665 1490.090 385.310 ;
        RECT 2503.630 383.090 2503.930 385.735 ;
        RECT 2903.830 383.090 2904.130 1084.775 ;
        RECT 1489.775 382.335 1490.105 382.665 ;
        RECT 1785.590 381.910 1786.770 383.090 ;
        RECT 1883.110 381.910 1884.290 383.090 ;
        RECT 1948.430 381.910 1949.610 383.090 ;
        RECT 2503.190 381.910 2504.370 383.090 ;
        RECT 2903.390 381.910 2904.570 383.090 ;
        RECT 1738.670 378.510 1739.850 379.690 ;
        RECT 1786.030 379.265 1786.330 381.910 ;
        RECT 1786.015 378.935 1786.345 379.265 ;
      LAYER met5 ;
        RECT 446.780 386.700 449.300 390.100 ;
        RECT 543.380 386.700 545.900 390.100 ;
        RECT 639.980 386.700 642.500 390.100 ;
        RECT 736.580 386.700 739.100 390.100 ;
        RECT 833.180 386.700 835.700 390.100 ;
        RECT 929.780 386.700 932.300 390.100 ;
        RECT 1026.380 386.700 1028.900 390.100 ;
        RECT 1122.980 386.700 1125.500 390.100 ;
        RECT 1219.580 386.700 1222.100 390.100 ;
        RECT 372.260 385.100 449.300 386.700 ;
        RECT 310.620 381.700 338.900 383.300 ;
        RECT 337.300 379.900 338.900 381.700 ;
        RECT 372.260 379.900 373.860 385.100 ;
        RECT 447.700 383.300 449.300 385.100 ;
        RECT 476.220 385.100 545.900 386.700 ;
        RECT 476.220 383.300 477.820 385.100 ;
        RECT 447.700 381.700 477.820 383.300 ;
        RECT 544.300 383.300 545.900 385.100 ;
        RECT 572.820 385.100 642.500 386.700 ;
        RECT 572.820 383.300 574.420 385.100 ;
        RECT 544.300 381.700 574.420 383.300 ;
        RECT 640.900 383.300 642.500 385.100 ;
        RECT 669.420 385.100 739.100 386.700 ;
        RECT 669.420 383.300 671.020 385.100 ;
        RECT 640.900 381.700 671.020 383.300 ;
        RECT 737.500 383.300 739.100 385.100 ;
        RECT 766.020 385.100 835.700 386.700 ;
        RECT 766.020 383.300 767.620 385.100 ;
        RECT 737.500 381.700 767.620 383.300 ;
        RECT 834.100 383.300 835.700 385.100 ;
        RECT 862.620 385.100 932.300 386.700 ;
        RECT 862.620 383.300 864.220 385.100 ;
        RECT 834.100 381.700 864.220 383.300 ;
        RECT 930.700 383.300 932.300 385.100 ;
        RECT 959.220 385.100 1028.900 386.700 ;
        RECT 959.220 383.300 960.820 385.100 ;
        RECT 930.700 381.700 960.820 383.300 ;
        RECT 1027.300 383.300 1028.900 385.100 ;
        RECT 1055.820 385.100 1125.500 386.700 ;
        RECT 1055.820 383.300 1057.420 385.100 ;
        RECT 1027.300 381.700 1057.420 383.300 ;
        RECT 1123.900 383.300 1125.500 385.100 ;
        RECT 1152.420 385.100 1222.100 386.700 ;
        RECT 1152.420 383.300 1154.020 385.100 ;
        RECT 1123.900 381.700 1154.020 383.300 ;
        RECT 1220.500 383.300 1222.100 385.100 ;
        RECT 1249.020 385.100 1316.860 386.700 ;
        RECT 1249.020 383.300 1250.620 385.100 ;
        RECT 1220.500 381.700 1250.620 383.300 ;
        RECT 337.300 378.300 373.860 379.900 ;
        RECT 1315.260 376.500 1316.860 385.100 ;
        RECT 1364.940 383.300 1367.460 390.100 ;
        RECT 1992.380 388.500 2046.420 390.100 ;
        RECT 1489.140 385.100 1498.100 386.700 ;
        RECT 1496.500 383.300 1498.100 385.100 ;
        RECT 1688.780 385.100 1705.100 386.700 ;
        RECT 1351.140 381.700 1407.940 383.300 ;
        RECT 1496.500 381.700 1545.940 383.300 ;
        RECT 1351.140 376.500 1352.740 381.700 ;
        RECT 1544.340 379.900 1545.940 381.700 ;
        RECT 1592.180 381.700 1607.580 383.300 ;
        RECT 1592.180 379.900 1593.780 381.700 ;
        RECT 1544.340 378.300 1593.780 379.900 ;
        RECT 1605.980 379.900 1607.580 381.700 ;
        RECT 1688.780 379.900 1690.380 385.100 ;
        RECT 1605.980 378.300 1690.380 379.900 ;
        RECT 1703.500 379.900 1705.100 385.100 ;
        RECT 1992.380 383.300 1993.980 388.500 ;
        RECT 2044.820 386.700 2046.420 388.500 ;
        RECT 2086.220 388.500 2091.500 390.100 ;
        RECT 2086.220 386.700 2087.820 388.500 ;
        RECT 2044.820 385.100 2087.820 386.700 ;
        RECT 1785.380 381.700 1800.780 383.300 ;
        RECT 1799.180 379.900 1800.780 381.700 ;
        RECT 1881.980 381.700 1885.280 383.300 ;
        RECT 1948.220 381.700 1993.980 383.300 ;
        RECT 2089.900 383.300 2091.500 388.500 ;
        RECT 2137.740 386.700 2140.260 390.100 ;
        RECT 2185.580 386.700 2188.100 390.100 ;
        RECT 2137.740 385.100 2188.100 386.700 ;
        RECT 2137.740 383.300 2139.340 385.100 ;
        RECT 2089.900 381.700 2139.340 383.300 ;
        RECT 2186.500 383.300 2188.100 385.100 ;
        RECT 2234.340 383.300 2236.860 390.100 ;
        RECT 2282.180 388.500 2381.300 390.100 ;
        RECT 2282.180 383.300 2283.780 388.500 ;
        RECT 2186.500 381.700 2283.780 383.300 ;
        RECT 2379.700 383.300 2381.300 388.500 ;
        RECT 2427.540 386.700 2430.060 390.100 ;
        RECT 2524.140 388.500 2529.420 390.100 ;
        RECT 2427.540 385.100 2475.140 386.700 ;
        RECT 2427.540 383.300 2429.140 385.100 ;
        RECT 2524.140 383.300 2525.740 388.500 ;
        RECT 2527.820 386.700 2529.420 388.500 ;
        RECT 2569.220 388.500 2574.500 390.100 ;
        RECT 2569.220 386.700 2570.820 388.500 ;
        RECT 2527.820 385.100 2570.820 386.700 ;
        RECT 2379.700 381.700 2429.140 383.300 ;
        RECT 2502.980 381.700 2525.740 383.300 ;
        RECT 2572.900 383.300 2574.500 388.500 ;
        RECT 2620.740 388.500 2673.860 390.100 ;
        RECT 2620.740 383.300 2622.340 388.500 ;
        RECT 2672.260 386.700 2673.860 388.500 ;
        RECT 2762.420 388.500 2767.700 390.100 ;
        RECT 2762.420 386.700 2764.020 388.500 ;
        RECT 2672.260 385.100 2764.020 386.700 ;
        RECT 2572.900 381.700 2622.340 383.300 ;
        RECT 2766.100 383.300 2767.700 388.500 ;
        RECT 2813.940 388.500 2836.700 390.100 ;
        RECT 2813.940 383.300 2815.540 388.500 ;
        RECT 2766.100 381.700 2815.540 383.300 ;
        RECT 2835.100 383.300 2836.700 388.500 ;
        RECT 2835.100 381.700 2904.780 383.300 ;
        RECT 1881.980 379.900 1883.580 381.700 ;
        RECT 1703.500 378.300 1740.060 379.900 ;
        RECT 1799.180 378.300 1883.580 379.900 ;
        RECT 1315.260 374.900 1352.740 376.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1150.990 1339.840 1151.310 1339.900 ;
        RECT 2898.990 1339.840 2899.310 1339.900 ;
        RECT 1150.990 1339.700 2899.310 1339.840 ;
        RECT 1150.990 1339.640 1151.310 1339.700 ;
        RECT 2898.990 1339.640 2899.310 1339.700 ;
      LAYER via ;
        RECT 1151.020 1339.640 1151.280 1339.900 ;
        RECT 2899.020 1339.640 2899.280 1339.900 ;
      LAYER met2 ;
        RECT 1151.020 1339.610 1151.280 1339.930 ;
        RECT 2899.020 1339.610 2899.280 1339.930 ;
        RECT 1151.080 1325.025 1151.220 1339.610 ;
        RECT 1150.970 1321.025 1151.250 1325.025 ;
        RECT 2899.080 1319.725 2899.220 1339.610 ;
        RECT 2899.010 1319.355 2899.290 1319.725 ;
      LAYER via2 ;
        RECT 2899.010 1319.400 2899.290 1319.680 ;
      LAYER met3 ;
        RECT 2898.985 1319.690 2899.315 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2898.985 1319.390 2924.800 1319.690 ;
        RECT 2898.985 1319.375 2899.315 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 305.970 1552.680 306.290 1552.740 ;
        RECT 2898.990 1552.680 2899.310 1552.740 ;
        RECT 305.970 1552.540 2899.310 1552.680 ;
        RECT 305.970 1552.480 306.290 1552.540 ;
        RECT 2898.990 1552.480 2899.310 1552.540 ;
      LAYER via ;
        RECT 306.000 1552.480 306.260 1552.740 ;
        RECT 2899.020 1552.480 2899.280 1552.740 ;
      LAYER met2 ;
        RECT 2899.010 1553.955 2899.290 1554.325 ;
        RECT 2899.080 1552.770 2899.220 1553.955 ;
        RECT 306.000 1552.450 306.260 1552.770 ;
        RECT 2899.020 1552.450 2899.280 1552.770 ;
        RECT 306.060 797.485 306.200 1552.450 ;
        RECT 305.990 797.115 306.270 797.485 ;
      LAYER via2 ;
        RECT 2899.010 1554.000 2899.290 1554.280 ;
        RECT 305.990 797.160 306.270 797.440 ;
      LAYER met3 ;
        RECT 2898.985 1554.290 2899.315 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2898.985 1553.990 2924.800 1554.290 ;
        RECT 2898.985 1553.975 2899.315 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 305.965 797.450 306.295 797.465 ;
        RECT 305.965 797.360 310.500 797.450 ;
        RECT 305.965 797.150 314.000 797.360 ;
        RECT 305.965 797.135 306.295 797.150 ;
        RECT 310.000 796.760 314.000 797.150 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1521.750 1787.280 1522.070 1787.340 ;
        RECT 2900.830 1787.280 2901.150 1787.340 ;
        RECT 1521.750 1787.140 2901.150 1787.280 ;
        RECT 1521.750 1787.080 1522.070 1787.140 ;
        RECT 2900.830 1787.080 2901.150 1787.140 ;
        RECT 1421.010 1255.860 1421.330 1255.920 ;
        RECT 1521.750 1255.860 1522.070 1255.920 ;
        RECT 1421.010 1255.720 1522.070 1255.860 ;
        RECT 1421.010 1255.660 1421.330 1255.720 ;
        RECT 1521.750 1255.660 1522.070 1255.720 ;
      LAYER via ;
        RECT 1521.780 1787.080 1522.040 1787.340 ;
        RECT 2900.860 1787.080 2901.120 1787.340 ;
        RECT 1421.040 1255.660 1421.300 1255.920 ;
        RECT 1521.780 1255.660 1522.040 1255.920 ;
      LAYER met2 ;
        RECT 2900.850 1789.235 2901.130 1789.605 ;
        RECT 2900.920 1787.370 2901.060 1789.235 ;
        RECT 1521.780 1787.050 1522.040 1787.370 ;
        RECT 2900.860 1787.050 2901.120 1787.370 ;
        RECT 1521.840 1255.950 1521.980 1787.050 ;
        RECT 1421.040 1255.630 1421.300 1255.950 ;
        RECT 1521.780 1255.630 1522.040 1255.950 ;
        RECT 1421.100 1250.365 1421.240 1255.630 ;
        RECT 1421.030 1249.995 1421.310 1250.365 ;
      LAYER via2 ;
        RECT 2900.850 1789.280 2901.130 1789.560 ;
        RECT 1421.030 1250.040 1421.310 1250.320 ;
      LAYER met3 ;
        RECT 2900.825 1789.570 2901.155 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.825 1789.270 2924.800 1789.570 ;
        RECT 2900.825 1789.255 2901.155 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 1421.005 1250.330 1421.335 1250.345 ;
        RECT 1408.060 1250.240 1421.335 1250.330 ;
        RECT 1404.305 1250.030 1421.335 1250.240 ;
        RECT 1404.305 1249.640 1408.305 1250.030 ;
        RECT 1421.005 1250.015 1421.335 1250.030 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1431.590 2021.880 1431.910 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 1431.590 2021.740 2901.150 2021.880 ;
        RECT 1431.590 2021.680 1431.910 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
        RECT 1000.110 214.440 1000.430 214.500 ;
        RECT 1431.590 214.440 1431.910 214.500 ;
        RECT 1000.110 214.300 1431.910 214.440 ;
        RECT 1000.110 214.240 1000.430 214.300 ;
        RECT 1431.590 214.240 1431.910 214.300 ;
      LAYER via ;
        RECT 1431.620 2021.680 1431.880 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
        RECT 1000.140 214.240 1000.400 214.500 ;
        RECT 1431.620 214.240 1431.880 214.500 ;
      LAYER met2 ;
        RECT 2900.850 2023.835 2901.130 2024.205 ;
        RECT 2900.920 2021.970 2901.060 2023.835 ;
        RECT 1431.620 2021.650 1431.880 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 1000.090 216.000 1000.370 220.000 ;
        RECT 1000.200 214.530 1000.340 216.000 ;
        RECT 1431.680 214.530 1431.820 2021.650 ;
        RECT 1000.140 214.210 1000.400 214.530 ;
        RECT 1431.620 214.210 1431.880 214.530 ;
      LAYER via2 ;
        RECT 2900.850 2023.880 2901.130 2024.160 ;
      LAYER met3 ;
        RECT 2900.825 2024.170 2901.155 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.825 2023.870 2924.800 2024.170 ;
        RECT 2900.825 2023.855 2901.155 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1497.000 2256.680 1499.440 2256.820 ;
        RECT 503.310 2256.480 503.630 2256.540 ;
        RECT 1497.000 2256.480 1497.140 2256.680 ;
        RECT 503.310 2256.340 1497.140 2256.480 ;
        RECT 1499.300 2256.480 1499.440 2256.680 ;
        RECT 2900.830 2256.480 2901.150 2256.540 ;
        RECT 1499.300 2256.340 2901.150 2256.480 ;
        RECT 503.310 2256.280 503.630 2256.340 ;
        RECT 2900.830 2256.280 2901.150 2256.340 ;
        RECT 497.790 1338.480 498.110 1338.540 ;
        RECT 503.310 1338.480 503.630 1338.540 ;
        RECT 497.790 1338.340 503.630 1338.480 ;
        RECT 497.790 1338.280 498.110 1338.340 ;
        RECT 503.310 1338.280 503.630 1338.340 ;
      LAYER via ;
        RECT 503.340 2256.280 503.600 2256.540 ;
        RECT 2900.860 2256.280 2901.120 2256.540 ;
        RECT 497.820 1338.280 498.080 1338.540 ;
        RECT 503.340 1338.280 503.600 1338.540 ;
      LAYER met2 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
        RECT 2900.920 2256.570 2901.060 2258.435 ;
        RECT 503.340 2256.250 503.600 2256.570 ;
        RECT 2900.860 2256.250 2901.120 2256.570 ;
        RECT 503.400 1338.570 503.540 2256.250 ;
        RECT 497.820 1338.250 498.080 1338.570 ;
        RECT 503.340 1338.250 503.600 1338.570 ;
        RECT 497.880 1325.025 498.020 1338.250 ;
        RECT 497.770 1321.025 498.050 1325.025 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
      LAYER met3 ;
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 760.395 1417.170 760.765 ;
        RECT 1416.960 634.965 1417.100 760.395 ;
        RECT 1416.890 634.595 1417.170 634.965 ;
        RECT 633.050 19.195 633.330 19.565 ;
        RECT 633.120 2.400 633.260 19.195 ;
        RECT 632.910 -4.800 633.470 2.400 ;
      LAYER via2 ;
        RECT 1416.890 760.440 1417.170 760.720 ;
        RECT 1416.890 634.640 1417.170 634.920 ;
        RECT 633.050 19.240 633.330 19.520 ;
      LAYER met3 ;
        RECT 1416.865 760.730 1417.195 760.745 ;
        RECT 1408.060 760.640 1417.195 760.730 ;
        RECT 1404.305 760.430 1417.195 760.640 ;
        RECT 1404.305 760.040 1408.305 760.430 ;
        RECT 1416.865 760.415 1417.195 760.430 ;
        RECT 1410.630 634.930 1411.010 634.940 ;
        RECT 1416.865 634.930 1417.195 634.945 ;
        RECT 1410.630 634.630 1417.195 634.930 ;
        RECT 1410.630 634.620 1411.010 634.630 ;
        RECT 1416.865 634.615 1417.195 634.630 ;
        RECT 633.025 19.530 633.355 19.545 ;
        RECT 1410.630 19.530 1411.010 19.540 ;
        RECT 633.025 19.230 1411.010 19.530 ;
        RECT 633.025 19.215 633.355 19.230 ;
        RECT 1410.630 19.220 1411.010 19.230 ;
      LAYER via3 ;
        RECT 1410.660 634.620 1410.980 634.940 ;
        RECT 1410.660 19.220 1410.980 19.540 ;
      LAYER met4 ;
        RECT 1410.655 634.615 1410.985 634.945 ;
        RECT 1410.670 19.545 1410.970 634.615 ;
        RECT 1410.655 19.215 1410.985 19.545 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1064.510 200.500 1064.830 200.560 ;
        RECT 1068.650 200.500 1068.970 200.560 ;
        RECT 1064.510 200.360 1068.970 200.500 ;
        RECT 1064.510 200.300 1064.830 200.360 ;
        RECT 1068.650 200.300 1068.970 200.360 ;
        RECT 1068.650 162.080 1068.970 162.140 ;
        RECT 2415.070 162.080 2415.390 162.140 ;
        RECT 1068.650 161.940 2415.390 162.080 ;
        RECT 1068.650 161.880 1068.970 161.940 ;
        RECT 2415.070 161.880 2415.390 161.940 ;
      LAYER via ;
        RECT 1064.540 200.300 1064.800 200.560 ;
        RECT 1068.680 200.300 1068.940 200.560 ;
        RECT 1068.680 161.880 1068.940 162.140 ;
        RECT 2415.100 161.880 2415.360 162.140 ;
      LAYER met2 ;
        RECT 1064.490 216.000 1064.770 220.000 ;
        RECT 1064.600 200.590 1064.740 216.000 ;
        RECT 1064.540 200.270 1064.800 200.590 ;
        RECT 1068.680 200.270 1068.940 200.590 ;
        RECT 1068.740 162.170 1068.880 200.270 ;
        RECT 1068.680 161.850 1068.940 162.170 ;
        RECT 2415.100 161.850 2415.360 162.170 ;
        RECT 2415.160 17.410 2415.300 161.850 ;
        RECT 2415.160 17.270 2417.600 17.410 ;
        RECT 2417.460 2.400 2417.600 17.270 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 710.075 286.950 710.445 ;
        RECT 286.740 17.525 286.880 710.075 ;
        RECT 286.670 17.155 286.950 17.525 ;
        RECT 2434.870 17.155 2435.150 17.525 ;
        RECT 2434.940 2.400 2435.080 17.155 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
      LAYER via2 ;
        RECT 286.670 710.120 286.950 710.400 ;
        RECT 286.670 17.200 286.950 17.480 ;
        RECT 2434.870 17.200 2435.150 17.480 ;
      LAYER met3 ;
        RECT 286.645 710.410 286.975 710.425 ;
        RECT 286.645 710.320 310.500 710.410 ;
        RECT 286.645 710.110 314.000 710.320 ;
        RECT 286.645 710.095 286.975 710.110 ;
        RECT 310.000 709.720 314.000 710.110 ;
        RECT 286.645 17.490 286.975 17.505 ;
        RECT 2434.845 17.490 2435.175 17.505 ;
        RECT 286.645 17.190 2435.175 17.490 ;
        RECT 286.645 17.175 286.975 17.190 ;
        RECT 2434.845 17.175 2435.175 17.190 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 280.670 1062.740 280.990 1062.800 ;
        RECT 296.770 1062.740 297.090 1062.800 ;
        RECT 280.670 1062.600 297.090 1062.740 ;
        RECT 280.670 1062.540 280.990 1062.600 ;
        RECT 296.770 1062.540 297.090 1062.600 ;
        RECT 1400.310 14.180 1400.630 14.240 ;
        RECT 2452.790 14.180 2453.110 14.240 ;
        RECT 1400.310 14.040 2453.110 14.180 ;
        RECT 1400.310 13.980 1400.630 14.040 ;
        RECT 2452.790 13.980 2453.110 14.040 ;
      LAYER via ;
        RECT 280.700 1062.540 280.960 1062.800 ;
        RECT 296.800 1062.540 297.060 1062.800 ;
        RECT 1400.340 13.980 1400.600 14.240 ;
        RECT 2452.820 13.980 2453.080 14.240 ;
      LAYER met2 ;
        RECT 296.790 1067.755 297.070 1068.125 ;
        RECT 296.860 1062.830 297.000 1067.755 ;
        RECT 280.700 1062.510 280.960 1062.830 ;
        RECT 296.800 1062.510 297.060 1062.830 ;
        RECT 280.760 20.245 280.900 1062.510 ;
        RECT 280.690 19.875 280.970 20.245 ;
        RECT 1400.330 19.875 1400.610 20.245 ;
        RECT 1400.400 14.270 1400.540 19.875 ;
        RECT 1400.340 13.950 1400.600 14.270 ;
        RECT 2452.820 13.950 2453.080 14.270 ;
        RECT 2452.880 2.400 2453.020 13.950 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
      LAYER via2 ;
        RECT 296.790 1067.800 297.070 1068.080 ;
        RECT 280.690 19.920 280.970 20.200 ;
        RECT 1400.330 19.920 1400.610 20.200 ;
      LAYER met3 ;
        RECT 296.765 1068.090 297.095 1068.105 ;
        RECT 296.765 1068.000 310.500 1068.090 ;
        RECT 296.765 1067.790 314.000 1068.000 ;
        RECT 296.765 1067.775 297.095 1067.790 ;
        RECT 310.000 1067.400 314.000 1067.790 ;
        RECT 280.665 20.210 280.995 20.225 ;
        RECT 1400.305 20.210 1400.635 20.225 ;
        RECT 280.665 19.910 1400.635 20.210 ;
        RECT 280.665 19.895 280.995 19.910 ;
        RECT 1400.305 19.895 1400.635 19.910 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.110 1336.780 448.430 1336.840 ;
        RECT 1352.470 1336.780 1352.790 1336.840 ;
        RECT 448.110 1336.640 1352.790 1336.780 ;
        RECT 448.110 1336.580 448.430 1336.640 ;
        RECT 1352.470 1336.580 1352.790 1336.640 ;
      LAYER via ;
        RECT 448.140 1336.580 448.400 1336.840 ;
        RECT 1352.500 1336.580 1352.760 1336.840 ;
      LAYER met2 ;
        RECT 448.140 1336.550 448.400 1336.870 ;
        RECT 1352.500 1336.550 1352.760 1336.870 ;
        RECT 448.200 1325.025 448.340 1336.550 ;
        RECT 1352.560 1333.325 1352.700 1336.550 ;
        RECT 1352.490 1332.955 1352.770 1333.325 ;
        RECT 2470.290 1332.955 2470.570 1333.325 ;
        RECT 448.090 1321.025 448.370 1325.025 ;
        RECT 2470.360 17.410 2470.500 1332.955 ;
        RECT 2470.360 17.270 2470.960 17.410 ;
        RECT 2470.820 2.400 2470.960 17.270 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
      LAYER via2 ;
        RECT 1352.490 1333.000 1352.770 1333.280 ;
        RECT 2470.290 1333.000 2470.570 1333.280 ;
      LAYER met3 ;
        RECT 1352.465 1333.290 1352.795 1333.305 ;
        RECT 2470.265 1333.290 2470.595 1333.305 ;
        RECT 1352.465 1332.990 2470.595 1333.290 ;
        RECT 1352.465 1332.975 1352.795 1332.990 ;
        RECT 2470.265 1332.975 2470.595 1332.990 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1131.760 1421.330 1131.820 ;
        RECT 2335.490 1131.760 2335.810 1131.820 ;
        RECT 1421.010 1131.620 2335.810 1131.760 ;
        RECT 1421.010 1131.560 1421.330 1131.620 ;
        RECT 2335.490 1131.560 2335.810 1131.620 ;
        RECT 2335.490 18.260 2335.810 18.320 ;
        RECT 2488.670 18.260 2488.990 18.320 ;
        RECT 2335.490 18.120 2488.990 18.260 ;
        RECT 2335.490 18.060 2335.810 18.120 ;
        RECT 2488.670 18.060 2488.990 18.120 ;
      LAYER via ;
        RECT 1421.040 1131.560 1421.300 1131.820 ;
        RECT 2335.520 1131.560 2335.780 1131.820 ;
        RECT 2335.520 18.060 2335.780 18.320 ;
        RECT 2488.700 18.060 2488.960 18.320 ;
      LAYER met2 ;
        RECT 1421.030 1133.035 1421.310 1133.405 ;
        RECT 1421.100 1131.850 1421.240 1133.035 ;
        RECT 1421.040 1131.530 1421.300 1131.850 ;
        RECT 2335.520 1131.530 2335.780 1131.850 ;
        RECT 2335.580 18.350 2335.720 1131.530 ;
        RECT 2335.520 18.030 2335.780 18.350 ;
        RECT 2488.700 18.030 2488.960 18.350 ;
        RECT 2488.760 2.400 2488.900 18.030 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1133.080 1421.310 1133.360 ;
      LAYER met3 ;
        RECT 1421.005 1133.370 1421.335 1133.385 ;
        RECT 1408.060 1133.280 1421.335 1133.370 ;
        RECT 1404.305 1133.070 1421.335 1133.280 ;
        RECT 1404.305 1132.680 1408.305 1133.070 ;
        RECT 1421.005 1133.055 1421.335 1133.070 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1202.510 201.180 1202.830 201.240 ;
        RECT 1206.190 201.180 1206.510 201.240 ;
        RECT 1202.510 201.040 1206.510 201.180 ;
        RECT 1202.510 200.980 1202.830 201.040 ;
        RECT 1206.190 200.980 1206.510 201.040 ;
        RECT 1206.190 128.080 1206.510 128.140 ;
        RECT 2504.770 128.080 2505.090 128.140 ;
        RECT 1206.190 127.940 2505.090 128.080 ;
        RECT 1206.190 127.880 1206.510 127.940 ;
        RECT 2504.770 127.880 2505.090 127.940 ;
      LAYER via ;
        RECT 1202.540 200.980 1202.800 201.240 ;
        RECT 1206.220 200.980 1206.480 201.240 ;
        RECT 1206.220 127.880 1206.480 128.140 ;
        RECT 2504.800 127.880 2505.060 128.140 ;
      LAYER met2 ;
        RECT 1202.490 216.000 1202.770 220.000 ;
        RECT 1202.600 201.270 1202.740 216.000 ;
        RECT 1202.540 200.950 1202.800 201.270 ;
        RECT 1206.220 200.950 1206.480 201.270 ;
        RECT 1206.280 128.170 1206.420 200.950 ;
        RECT 1206.220 127.850 1206.480 128.170 ;
        RECT 2504.800 127.850 2505.060 128.170 ;
        RECT 2504.860 17.410 2505.000 127.850 ;
        RECT 2504.860 17.270 2506.380 17.410 ;
        RECT 2506.240 2.400 2506.380 17.270 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 287.110 713.220 287.430 713.280 ;
        RECT 296.770 713.220 297.090 713.280 ;
        RECT 287.110 713.080 297.090 713.220 ;
        RECT 287.110 713.020 287.430 713.080 ;
        RECT 296.770 713.020 297.090 713.080 ;
      LAYER via ;
        RECT 287.140 713.020 287.400 713.280 ;
        RECT 296.800 713.020 297.060 713.280 ;
      LAYER met2 ;
        RECT 296.790 716.875 297.070 717.245 ;
        RECT 296.860 713.310 297.000 716.875 ;
        RECT 287.140 712.990 287.400 713.310 ;
        RECT 296.800 712.990 297.060 713.310 ;
        RECT 287.200 16.845 287.340 712.990 ;
        RECT 287.130 16.475 287.410 16.845 ;
        RECT 2524.110 16.475 2524.390 16.845 ;
        RECT 2524.180 2.400 2524.320 16.475 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
      LAYER via2 ;
        RECT 296.790 716.920 297.070 717.200 ;
        RECT 287.130 16.520 287.410 16.800 ;
        RECT 2524.110 16.520 2524.390 16.800 ;
      LAYER met3 ;
        RECT 296.765 717.210 297.095 717.225 ;
        RECT 296.765 717.120 310.500 717.210 ;
        RECT 296.765 716.910 314.000 717.120 ;
        RECT 296.765 716.895 297.095 716.910 ;
        RECT 310.000 716.520 314.000 716.910 ;
        RECT 287.105 16.810 287.435 16.825 ;
        RECT 2524.085 16.810 2524.415 16.825 ;
        RECT 287.105 16.510 2524.415 16.810 ;
        RECT 287.105 16.495 287.435 16.510 ;
        RECT 2524.085 16.495 2524.415 16.510 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1166.440 1421.330 1166.500 ;
        RECT 1541.990 1166.440 1542.310 1166.500 ;
        RECT 1421.010 1166.300 1542.310 1166.440 ;
        RECT 1421.010 1166.240 1421.330 1166.300 ;
        RECT 1541.990 1166.240 1542.310 1166.300 ;
        RECT 1541.990 59.060 1542.310 59.120 ;
        RECT 2539.270 59.060 2539.590 59.120 ;
        RECT 1541.990 58.920 2539.590 59.060 ;
        RECT 1541.990 58.860 1542.310 58.920 ;
        RECT 2539.270 58.860 2539.590 58.920 ;
      LAYER via ;
        RECT 1421.040 1166.240 1421.300 1166.500 ;
        RECT 1542.020 1166.240 1542.280 1166.500 ;
        RECT 1542.020 58.860 1542.280 59.120 ;
        RECT 2539.300 58.860 2539.560 59.120 ;
      LAYER met2 ;
        RECT 1421.030 1169.755 1421.310 1170.125 ;
        RECT 1421.100 1166.530 1421.240 1169.755 ;
        RECT 1421.040 1166.210 1421.300 1166.530 ;
        RECT 1542.020 1166.210 1542.280 1166.530 ;
        RECT 1542.080 59.150 1542.220 1166.210 ;
        RECT 1542.020 58.830 1542.280 59.150 ;
        RECT 2539.300 58.830 2539.560 59.150 ;
        RECT 2539.360 17.410 2539.500 58.830 ;
        RECT 2539.360 17.270 2542.260 17.410 ;
        RECT 2542.120 2.400 2542.260 17.270 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1169.800 1421.310 1170.080 ;
      LAYER met3 ;
        RECT 1421.005 1170.090 1421.335 1170.105 ;
        RECT 1408.060 1170.000 1421.335 1170.090 ;
        RECT 1404.305 1169.790 1421.335 1170.000 ;
        RECT 1404.305 1169.400 1408.305 1169.790 ;
        RECT 1421.005 1169.775 1421.335 1169.790 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 1326.835 325.130 1327.205 ;
        RECT 2559.990 1326.835 2560.270 1327.205 ;
        RECT 324.920 1325.025 325.060 1326.835 ;
        RECT 324.810 1321.025 325.090 1325.025 ;
        RECT 2560.060 2.400 2560.200 1326.835 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
      LAYER via2 ;
        RECT 324.850 1326.880 325.130 1327.160 ;
        RECT 2559.990 1326.880 2560.270 1327.160 ;
      LAYER met3 ;
        RECT 324.825 1327.170 325.155 1327.185 ;
        RECT 2559.965 1327.170 2560.295 1327.185 ;
        RECT 324.825 1326.870 2560.295 1327.170 ;
        RECT 324.825 1326.855 325.155 1326.870 ;
        RECT 2559.965 1326.855 2560.295 1326.870 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 871.310 200.500 871.630 200.560 ;
        RECT 875.910 200.500 876.230 200.560 ;
        RECT 871.310 200.360 876.230 200.500 ;
        RECT 871.310 200.300 871.630 200.360 ;
        RECT 875.910 200.300 876.230 200.360 ;
        RECT 875.910 93.400 876.230 93.460 ;
        RECT 2573.770 93.400 2574.090 93.460 ;
        RECT 875.910 93.260 2574.090 93.400 ;
        RECT 875.910 93.200 876.230 93.260 ;
        RECT 2573.770 93.200 2574.090 93.260 ;
      LAYER via ;
        RECT 871.340 200.300 871.600 200.560 ;
        RECT 875.940 200.300 876.200 200.560 ;
        RECT 875.940 93.200 876.200 93.460 ;
        RECT 2573.800 93.200 2574.060 93.460 ;
      LAYER met2 ;
        RECT 871.290 216.000 871.570 220.000 ;
        RECT 871.400 200.590 871.540 216.000 ;
        RECT 871.340 200.270 871.600 200.590 ;
        RECT 875.940 200.270 876.200 200.590 ;
        RECT 876.000 93.490 876.140 200.270 ;
        RECT 875.940 93.170 876.200 93.490 ;
        RECT 2573.800 93.170 2574.060 93.490 ;
        RECT 2573.860 17.410 2574.000 93.170 ;
        RECT 2573.860 17.270 2578.140 17.410 ;
        RECT 2578.000 2.400 2578.140 17.270 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 813.350 107.340 813.670 107.400 ;
        RECT 1411.350 107.340 1411.670 107.400 ;
        RECT 813.350 107.200 1411.670 107.340 ;
        RECT 813.350 107.140 813.670 107.200 ;
        RECT 1411.350 107.140 1411.670 107.200 ;
      LAYER via ;
        RECT 813.380 107.140 813.640 107.400 ;
        RECT 1411.380 107.140 1411.640 107.400 ;
      LAYER met2 ;
        RECT 1411.370 255.835 1411.650 256.205 ;
        RECT 1411.440 107.430 1411.580 255.835 ;
        RECT 813.380 107.110 813.640 107.430 ;
        RECT 1411.380 107.110 1411.640 107.430 ;
        RECT 813.440 17.410 813.580 107.110 ;
        RECT 811.600 17.270 813.580 17.410 ;
        RECT 811.600 2.400 811.740 17.270 ;
        RECT 811.390 -4.800 811.950 2.400 ;
      LAYER via2 ;
        RECT 1411.370 255.880 1411.650 256.160 ;
      LAYER met3 ;
        RECT 1411.345 256.170 1411.675 256.185 ;
        RECT 1408.060 256.080 1411.675 256.170 ;
        RECT 1404.305 255.870 1411.675 256.080 ;
        RECT 1404.305 255.480 1408.305 255.870 ;
        RECT 1411.345 255.855 1411.675 255.870 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 843.710 1340.180 844.030 1340.240 ;
        RECT 2594.470 1340.180 2594.790 1340.240 ;
        RECT 843.710 1340.040 2594.790 1340.180 ;
        RECT 843.710 1339.980 844.030 1340.040 ;
        RECT 2594.470 1339.980 2594.790 1340.040 ;
      LAYER via ;
        RECT 843.740 1339.980 844.000 1340.240 ;
        RECT 2594.500 1339.980 2594.760 1340.240 ;
      LAYER met2 ;
        RECT 843.740 1339.950 844.000 1340.270 ;
        RECT 2594.500 1339.950 2594.760 1340.270 ;
        RECT 843.800 1325.025 843.940 1339.950 ;
        RECT 843.690 1321.025 843.970 1325.025 ;
        RECT 2594.560 17.410 2594.700 1339.950 ;
        RECT 2594.560 17.270 2595.620 17.410 ;
        RECT 2595.480 2.400 2595.620 17.270 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.030 1339.160 725.350 1339.220 ;
        RECT 2608.270 1339.160 2608.590 1339.220 ;
        RECT 725.030 1339.020 2608.590 1339.160 ;
        RECT 725.030 1338.960 725.350 1339.020 ;
        RECT 2608.270 1338.960 2608.590 1339.020 ;
      LAYER via ;
        RECT 725.060 1338.960 725.320 1339.220 ;
        RECT 2608.300 1338.960 2608.560 1339.220 ;
      LAYER met2 ;
        RECT 725.060 1338.930 725.320 1339.250 ;
        RECT 2608.300 1338.930 2608.560 1339.250 ;
        RECT 725.120 1325.025 725.260 1338.930 ;
        RECT 725.010 1321.025 725.290 1325.025 ;
        RECT 2608.360 17.410 2608.500 1338.930 ;
        RECT 2608.360 17.270 2613.560 17.410 ;
        RECT 2613.420 2.400 2613.560 17.270 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 279.290 372.880 279.610 372.940 ;
        RECT 296.770 372.880 297.090 372.940 ;
        RECT 279.290 372.740 297.090 372.880 ;
        RECT 279.290 372.680 279.610 372.740 ;
        RECT 296.770 372.680 297.090 372.740 ;
      LAYER via ;
        RECT 279.320 372.680 279.580 372.940 ;
        RECT 296.800 372.680 297.060 372.940 ;
      LAYER met2 ;
        RECT 279.320 372.650 279.580 372.970 ;
        RECT 296.790 372.795 297.070 373.165 ;
        RECT 296.800 372.650 297.060 372.795 ;
        RECT 279.380 33.845 279.520 372.650 ;
        RECT 279.310 33.475 279.590 33.845 ;
        RECT 2631.290 33.475 2631.570 33.845 ;
        RECT 2631.360 2.400 2631.500 33.475 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
      LAYER via2 ;
        RECT 296.790 372.840 297.070 373.120 ;
        RECT 279.310 33.520 279.590 33.800 ;
        RECT 2631.290 33.520 2631.570 33.800 ;
      LAYER met3 ;
        RECT 296.765 373.130 297.095 373.145 ;
        RECT 296.765 373.040 310.500 373.130 ;
        RECT 296.765 372.830 314.000 373.040 ;
        RECT 296.765 372.815 297.095 372.830 ;
        RECT 310.000 372.440 314.000 372.830 ;
        RECT 279.285 33.810 279.615 33.825 ;
        RECT 2631.265 33.810 2631.595 33.825 ;
        RECT 279.285 33.510 2631.595 33.810 ;
        RECT 279.285 33.495 279.615 33.510 ;
        RECT 2631.265 33.495 2631.595 33.510 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1415.950 1304.480 1416.270 1304.540 ;
        RECT 1521.290 1304.480 1521.610 1304.540 ;
        RECT 1415.950 1304.340 1521.610 1304.480 ;
        RECT 1415.950 1304.280 1416.270 1304.340 ;
        RECT 1521.290 1304.280 1521.610 1304.340 ;
        RECT 1521.290 80.480 1521.610 80.540 ;
        RECT 2643.230 80.480 2643.550 80.540 ;
        RECT 1521.290 80.340 2643.550 80.480 ;
        RECT 1521.290 80.280 1521.610 80.340 ;
        RECT 2643.230 80.280 2643.550 80.340 ;
        RECT 2643.230 18.260 2643.550 18.320 ;
        RECT 2649.210 18.260 2649.530 18.320 ;
        RECT 2643.230 18.120 2649.530 18.260 ;
        RECT 2643.230 18.060 2643.550 18.120 ;
        RECT 2649.210 18.060 2649.530 18.120 ;
      LAYER via ;
        RECT 1415.980 1304.280 1416.240 1304.540 ;
        RECT 1521.320 1304.280 1521.580 1304.540 ;
        RECT 1521.320 80.280 1521.580 80.540 ;
        RECT 2643.260 80.280 2643.520 80.540 ;
        RECT 2643.260 18.060 2643.520 18.320 ;
        RECT 2649.240 18.060 2649.500 18.320 ;
      LAYER met2 ;
        RECT 1415.970 1308.475 1416.250 1308.845 ;
        RECT 1416.040 1304.570 1416.180 1308.475 ;
        RECT 1415.980 1304.250 1416.240 1304.570 ;
        RECT 1521.320 1304.250 1521.580 1304.570 ;
        RECT 1521.380 80.570 1521.520 1304.250 ;
        RECT 1521.320 80.250 1521.580 80.570 ;
        RECT 2643.260 80.250 2643.520 80.570 ;
        RECT 2643.320 18.350 2643.460 80.250 ;
        RECT 2643.260 18.030 2643.520 18.350 ;
        RECT 2649.240 18.030 2649.500 18.350 ;
        RECT 2649.300 2.400 2649.440 18.030 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
      LAYER via2 ;
        RECT 1415.970 1308.520 1416.250 1308.800 ;
      LAYER met3 ;
        RECT 1415.945 1308.810 1416.275 1308.825 ;
        RECT 1408.060 1308.720 1416.275 1308.810 ;
        RECT 1404.305 1308.510 1416.275 1308.720 ;
        RECT 1404.305 1308.120 1408.305 1308.510 ;
        RECT 1415.945 1308.495 1416.275 1308.510 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1014.830 200.500 1015.150 200.560 ;
        RECT 1020.350 200.500 1020.670 200.560 ;
        RECT 1014.830 200.360 1020.670 200.500 ;
        RECT 1014.830 200.300 1015.150 200.360 ;
        RECT 1020.350 200.300 1020.670 200.360 ;
        RECT 1020.350 87.280 1020.670 87.340 ;
        RECT 2663.470 87.280 2663.790 87.340 ;
        RECT 1020.350 87.140 2663.790 87.280 ;
        RECT 1020.350 87.080 1020.670 87.140 ;
        RECT 2663.470 87.080 2663.790 87.140 ;
      LAYER via ;
        RECT 1014.860 200.300 1015.120 200.560 ;
        RECT 1020.380 200.300 1020.640 200.560 ;
        RECT 1020.380 87.080 1020.640 87.340 ;
        RECT 2663.500 87.080 2663.760 87.340 ;
      LAYER met2 ;
        RECT 1014.810 216.000 1015.090 220.000 ;
        RECT 1014.920 200.590 1015.060 216.000 ;
        RECT 1014.860 200.270 1015.120 200.590 ;
        RECT 1020.380 200.270 1020.640 200.590 ;
        RECT 1020.440 87.370 1020.580 200.270 ;
        RECT 1020.380 87.050 1020.640 87.370 ;
        RECT 2663.500 87.050 2663.760 87.370 ;
        RECT 2663.560 17.410 2663.700 87.050 ;
        RECT 2663.560 17.270 2667.380 17.410 ;
        RECT 2667.240 2.400 2667.380 17.270 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 1334.315 537.650 1334.685 ;
        RECT 537.440 1325.025 537.580 1334.315 ;
        RECT 537.330 1321.025 537.610 1325.025 ;
        RECT 2684.650 17.155 2684.930 17.525 ;
        RECT 2684.720 2.400 2684.860 17.155 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
      LAYER via2 ;
        RECT 537.370 1334.360 537.650 1334.640 ;
        RECT 2684.650 17.200 2684.930 17.480 ;
      LAYER met3 ;
        RECT 1400.510 1338.050 1400.890 1338.060 ;
        RECT 1448.350 1338.050 1448.730 1338.060 ;
        RECT 1400.510 1337.750 1448.730 1338.050 ;
        RECT 1400.510 1337.740 1400.890 1337.750 ;
        RECT 1448.350 1337.740 1448.730 1337.750 ;
        RECT 1460.310 1338.050 1460.690 1338.060 ;
        RECT 1473.190 1338.050 1473.570 1338.060 ;
        RECT 1460.310 1337.750 1473.570 1338.050 ;
        RECT 1460.310 1337.740 1460.690 1337.750 ;
        RECT 1473.190 1337.740 1473.570 1337.750 ;
        RECT 1207.310 1336.690 1207.690 1336.700 ;
        RECT 1222.950 1336.690 1223.330 1336.700 ;
        RECT 1207.310 1336.390 1223.330 1336.690 ;
        RECT 1207.310 1336.380 1207.690 1336.390 ;
        RECT 1222.950 1336.380 1223.330 1336.390 ;
        RECT 537.345 1334.660 537.675 1334.665 ;
        RECT 537.345 1334.650 537.930 1334.660 ;
        RECT 537.120 1334.350 537.930 1334.650 ;
        RECT 537.345 1334.340 537.930 1334.350 ;
        RECT 1497.110 1334.650 1497.490 1334.660 ;
        RECT 1544.950 1334.650 1545.330 1334.660 ;
        RECT 1497.110 1334.350 1545.330 1334.650 ;
        RECT 1497.110 1334.340 1497.490 1334.350 ;
        RECT 1544.950 1334.340 1545.330 1334.350 ;
        RECT 1604.750 1334.650 1605.130 1334.660 ;
        RECT 1641.550 1334.650 1641.930 1334.660 ;
        RECT 1604.750 1334.350 1641.930 1334.650 ;
        RECT 1604.750 1334.340 1605.130 1334.350 ;
        RECT 1641.550 1334.340 1641.930 1334.350 ;
        RECT 1690.310 1334.650 1690.690 1334.660 ;
        RECT 1738.150 1334.650 1738.530 1334.660 ;
        RECT 1690.310 1334.350 1738.530 1334.650 ;
        RECT 1690.310 1334.340 1690.690 1334.350 ;
        RECT 1738.150 1334.340 1738.530 1334.350 ;
        RECT 1786.910 1334.650 1787.290 1334.660 ;
        RECT 1834.750 1334.650 1835.130 1334.660 ;
        RECT 1786.910 1334.350 1835.130 1334.650 ;
        RECT 1786.910 1334.340 1787.290 1334.350 ;
        RECT 1834.750 1334.340 1835.130 1334.350 ;
        RECT 1884.430 1334.650 1884.810 1334.660 ;
        RECT 1931.350 1334.650 1931.730 1334.660 ;
        RECT 1884.430 1334.350 1931.730 1334.650 ;
        RECT 1884.430 1334.340 1884.810 1334.350 ;
        RECT 1931.350 1334.340 1931.730 1334.350 ;
        RECT 1980.110 1334.650 1980.490 1334.660 ;
        RECT 2027.950 1334.650 2028.330 1334.660 ;
        RECT 1980.110 1334.350 2028.330 1334.650 ;
        RECT 1980.110 1334.340 1980.490 1334.350 ;
        RECT 2027.950 1334.340 2028.330 1334.350 ;
        RECT 2087.750 1334.650 2088.130 1334.660 ;
        RECT 2124.550 1334.650 2124.930 1334.660 ;
        RECT 2087.750 1334.350 2124.930 1334.650 ;
        RECT 2087.750 1334.340 2088.130 1334.350 ;
        RECT 2124.550 1334.340 2124.930 1334.350 ;
        RECT 2184.350 1334.650 2184.730 1334.660 ;
        RECT 2221.150 1334.650 2221.530 1334.660 ;
        RECT 2184.350 1334.350 2221.530 1334.650 ;
        RECT 2184.350 1334.340 2184.730 1334.350 ;
        RECT 2221.150 1334.340 2221.530 1334.350 ;
        RECT 2280.950 1334.650 2281.330 1334.660 ;
        RECT 2317.750 1334.650 2318.130 1334.660 ;
        RECT 2280.950 1334.350 2318.130 1334.650 ;
        RECT 2280.950 1334.340 2281.330 1334.350 ;
        RECT 2317.750 1334.340 2318.130 1334.350 ;
        RECT 2377.550 1334.650 2377.930 1334.660 ;
        RECT 2414.350 1334.650 2414.730 1334.660 ;
        RECT 2377.550 1334.350 2414.730 1334.650 ;
        RECT 2377.550 1334.340 2377.930 1334.350 ;
        RECT 2414.350 1334.340 2414.730 1334.350 ;
        RECT 2464.030 1334.650 2464.410 1334.660 ;
        RECT 2510.950 1334.650 2511.330 1334.660 ;
        RECT 2464.030 1334.350 2511.330 1334.650 ;
        RECT 2464.030 1334.340 2464.410 1334.350 ;
        RECT 2510.950 1334.340 2511.330 1334.350 ;
        RECT 2559.710 1334.650 2560.090 1334.660 ;
        RECT 2607.550 1334.650 2607.930 1334.660 ;
        RECT 2559.710 1334.350 2607.930 1334.650 ;
        RECT 2559.710 1334.340 2560.090 1334.350 ;
        RECT 2607.550 1334.340 2607.930 1334.350 ;
        RECT 2669.190 1334.650 2669.570 1334.660 ;
        RECT 2683.910 1334.650 2684.290 1334.660 ;
        RECT 2669.190 1334.350 2684.290 1334.650 ;
        RECT 2669.190 1334.340 2669.570 1334.350 ;
        RECT 2683.910 1334.340 2684.290 1334.350 ;
        RECT 537.345 1334.335 537.675 1334.340 ;
        RECT 1159.470 1331.250 1159.850 1331.260 ;
        RECT 1206.390 1331.250 1206.770 1331.260 ;
        RECT 1159.470 1330.950 1206.770 1331.250 ;
        RECT 1159.470 1330.940 1159.850 1330.950 ;
        RECT 1206.390 1330.940 1206.770 1330.950 ;
        RECT 2683.910 17.490 2684.290 17.500 ;
        RECT 2684.625 17.490 2684.955 17.505 ;
        RECT 2683.910 17.190 2684.955 17.490 ;
        RECT 2683.910 17.180 2684.290 17.190 ;
        RECT 2684.625 17.175 2684.955 17.190 ;
      LAYER via3 ;
        RECT 1400.540 1337.740 1400.860 1338.060 ;
        RECT 1448.380 1337.740 1448.700 1338.060 ;
        RECT 1460.340 1337.740 1460.660 1338.060 ;
        RECT 1473.220 1337.740 1473.540 1338.060 ;
        RECT 1207.340 1336.380 1207.660 1336.700 ;
        RECT 1222.980 1336.380 1223.300 1336.700 ;
        RECT 537.580 1334.340 537.900 1334.660 ;
        RECT 1497.140 1334.340 1497.460 1334.660 ;
        RECT 1544.980 1334.340 1545.300 1334.660 ;
        RECT 1604.780 1334.340 1605.100 1334.660 ;
        RECT 1641.580 1334.340 1641.900 1334.660 ;
        RECT 1690.340 1334.340 1690.660 1334.660 ;
        RECT 1738.180 1334.340 1738.500 1334.660 ;
        RECT 1786.940 1334.340 1787.260 1334.660 ;
        RECT 1834.780 1334.340 1835.100 1334.660 ;
        RECT 1884.460 1334.340 1884.780 1334.660 ;
        RECT 1931.380 1334.340 1931.700 1334.660 ;
        RECT 1980.140 1334.340 1980.460 1334.660 ;
        RECT 2027.980 1334.340 2028.300 1334.660 ;
        RECT 2087.780 1334.340 2088.100 1334.660 ;
        RECT 2124.580 1334.340 2124.900 1334.660 ;
        RECT 2184.380 1334.340 2184.700 1334.660 ;
        RECT 2221.180 1334.340 2221.500 1334.660 ;
        RECT 2280.980 1334.340 2281.300 1334.660 ;
        RECT 2317.780 1334.340 2318.100 1334.660 ;
        RECT 2377.580 1334.340 2377.900 1334.660 ;
        RECT 2414.380 1334.340 2414.700 1334.660 ;
        RECT 2464.060 1334.340 2464.380 1334.660 ;
        RECT 2510.980 1334.340 2511.300 1334.660 ;
        RECT 2559.740 1334.340 2560.060 1334.660 ;
        RECT 2607.580 1334.340 2607.900 1334.660 ;
        RECT 2669.220 1334.340 2669.540 1334.660 ;
        RECT 2683.940 1334.340 2684.260 1334.660 ;
        RECT 1159.500 1330.940 1159.820 1331.260 ;
        RECT 1206.420 1330.940 1206.740 1331.260 ;
        RECT 2683.940 17.180 2684.260 17.500 ;
      LAYER met4 ;
        RECT 1400.535 1337.735 1400.865 1338.065 ;
        RECT 1207.335 1336.375 1207.665 1336.705 ;
        RECT 1222.975 1336.375 1223.305 1336.705 ;
        RECT 1207.350 1335.090 1207.650 1336.375 ;
        RECT 1222.990 1335.090 1223.290 1336.375 ;
        RECT 1400.550 1335.090 1400.850 1337.735 ;
        RECT 1447.950 1337.310 1449.130 1338.490 ;
        RECT 1459.910 1337.310 1461.090 1338.490 ;
        RECT 1473.215 1337.735 1473.545 1338.065 ;
        RECT 1473.230 1335.090 1473.530 1337.735 ;
        RECT 2668.790 1337.310 2669.970 1338.490 ;
        RECT 537.150 1333.910 538.330 1335.090 ;
        RECT 1159.070 1333.910 1160.250 1335.090 ;
        RECT 1206.910 1333.910 1208.090 1335.090 ;
        RECT 1222.550 1333.910 1223.730 1335.090 ;
        RECT 1400.110 1333.910 1401.290 1335.090 ;
        RECT 1472.790 1333.910 1473.970 1335.090 ;
        RECT 1496.710 1333.910 1497.890 1335.090 ;
        RECT 1544.975 1334.335 1545.305 1334.665 ;
        RECT 1159.510 1331.265 1159.810 1333.910 ;
        RECT 1544.990 1331.690 1545.290 1334.335 ;
        RECT 1604.350 1333.910 1605.530 1335.090 ;
        RECT 1641.575 1334.335 1641.905 1334.665 ;
        RECT 1641.590 1331.690 1641.890 1334.335 ;
        RECT 1689.910 1333.910 1691.090 1335.090 ;
        RECT 1738.175 1334.335 1738.505 1334.665 ;
        RECT 1738.190 1331.690 1738.490 1334.335 ;
        RECT 1786.510 1333.910 1787.690 1335.090 ;
        RECT 1834.775 1334.335 1835.105 1334.665 ;
        RECT 1834.790 1331.690 1835.090 1334.335 ;
        RECT 1884.030 1333.910 1885.210 1335.090 ;
        RECT 1931.375 1334.335 1931.705 1334.665 ;
        RECT 1931.390 1331.690 1931.690 1334.335 ;
        RECT 1979.710 1333.910 1980.890 1335.090 ;
        RECT 2027.975 1334.335 2028.305 1334.665 ;
        RECT 2027.990 1331.690 2028.290 1334.335 ;
        RECT 2087.350 1333.910 2088.530 1335.090 ;
        RECT 2124.575 1334.335 2124.905 1334.665 ;
        RECT 2124.590 1331.690 2124.890 1334.335 ;
        RECT 2183.950 1333.910 2185.130 1335.090 ;
        RECT 2221.175 1334.335 2221.505 1334.665 ;
        RECT 2221.190 1331.690 2221.490 1334.335 ;
        RECT 2280.550 1333.910 2281.730 1335.090 ;
        RECT 2317.775 1334.335 2318.105 1334.665 ;
        RECT 2317.790 1331.690 2318.090 1334.335 ;
        RECT 2377.150 1333.910 2378.330 1335.090 ;
        RECT 2414.375 1334.335 2414.705 1334.665 ;
        RECT 2414.390 1331.690 2414.690 1334.335 ;
        RECT 2463.630 1333.910 2464.810 1335.090 ;
        RECT 2510.975 1334.335 2511.305 1334.665 ;
        RECT 2510.990 1331.690 2511.290 1334.335 ;
        RECT 2559.310 1333.910 2560.490 1335.090 ;
        RECT 2669.230 1334.665 2669.530 1337.310 ;
        RECT 2607.575 1334.335 2607.905 1334.665 ;
        RECT 2669.215 1334.335 2669.545 1334.665 ;
        RECT 2683.935 1334.335 2684.265 1334.665 ;
        RECT 2607.590 1331.690 2607.890 1334.335 ;
        RECT 1159.495 1330.935 1159.825 1331.265 ;
        RECT 1205.990 1330.510 1207.170 1331.690 ;
        RECT 1544.550 1330.510 1545.730 1331.690 ;
        RECT 1641.150 1330.510 1642.330 1331.690 ;
        RECT 1737.750 1330.510 1738.930 1331.690 ;
        RECT 1834.350 1330.510 1835.530 1331.690 ;
        RECT 1930.950 1330.510 1932.130 1331.690 ;
        RECT 2027.550 1330.510 2028.730 1331.690 ;
        RECT 2124.150 1330.510 2125.330 1331.690 ;
        RECT 2220.750 1330.510 2221.930 1331.690 ;
        RECT 2317.350 1330.510 2318.530 1331.690 ;
        RECT 2413.950 1330.510 2415.130 1331.690 ;
        RECT 2510.550 1330.510 2511.730 1331.690 ;
        RECT 2607.150 1330.510 2608.330 1331.690 ;
        RECT 2683.950 17.505 2684.250 1334.335 ;
        RECT 2683.935 17.175 2684.265 17.505 ;
      LAYER met5 ;
        RECT 545.220 1337.100 594.660 1338.700 ;
        RECT 545.220 1335.300 546.820 1337.100 ;
        RECT 536.940 1333.700 546.820 1335.300 ;
        RECT 593.060 1335.300 594.660 1337.100 ;
        RECT 662.060 1337.100 712.420 1338.700 ;
        RECT 662.060 1335.300 663.660 1337.100 ;
        RECT 593.060 1333.700 663.660 1335.300 ;
        RECT 710.820 1335.300 712.420 1337.100 ;
        RECT 758.660 1337.100 809.020 1338.700 ;
        RECT 758.660 1335.300 760.260 1337.100 ;
        RECT 710.820 1333.700 760.260 1335.300 ;
        RECT 807.420 1335.300 809.020 1337.100 ;
        RECT 855.260 1337.100 905.620 1338.700 ;
        RECT 855.260 1335.300 856.860 1337.100 ;
        RECT 807.420 1333.700 856.860 1335.300 ;
        RECT 904.020 1335.300 905.620 1337.100 ;
        RECT 951.860 1337.100 1001.300 1338.700 ;
        RECT 951.860 1335.300 953.460 1337.100 ;
        RECT 904.020 1333.700 953.460 1335.300 ;
        RECT 999.700 1335.300 1001.300 1337.100 ;
        RECT 1028.220 1337.100 1126.420 1338.700 ;
        RECT 1028.220 1335.300 1029.820 1337.100 ;
        RECT 999.700 1333.700 1029.820 1335.300 ;
        RECT 1124.820 1335.300 1126.420 1337.100 ;
        RECT 1269.260 1337.100 1304.900 1338.700 ;
        RECT 1447.740 1337.100 1461.300 1338.700 ;
        RECT 2621.660 1337.100 2670.180 1338.700 ;
        RECT 1269.260 1335.300 1270.860 1337.100 ;
        RECT 1124.820 1333.700 1160.460 1335.300 ;
        RECT 1206.700 1331.900 1208.300 1335.300 ;
        RECT 1222.340 1333.700 1270.860 1335.300 ;
        RECT 1303.300 1335.300 1304.900 1337.100 ;
        RECT 1303.300 1333.700 1401.500 1335.300 ;
        RECT 1472.580 1333.700 1498.100 1335.300 ;
        RECT 1559.060 1333.700 1605.740 1335.300 ;
        RECT 1655.660 1333.700 1691.300 1335.300 ;
        RECT 1752.260 1333.700 1787.900 1335.300 ;
        RECT 1848.860 1333.700 1885.420 1335.300 ;
        RECT 1945.460 1333.700 1981.100 1335.300 ;
        RECT 2042.060 1333.700 2088.740 1335.300 ;
        RECT 2138.660 1333.700 2185.340 1335.300 ;
        RECT 2235.260 1333.700 2281.940 1335.300 ;
        RECT 2331.860 1333.700 2378.540 1335.300 ;
        RECT 2428.460 1333.700 2465.020 1335.300 ;
        RECT 2525.060 1333.700 2560.700 1335.300 ;
        RECT 1559.060 1331.900 1560.660 1333.700 ;
        RECT 1655.660 1331.900 1657.260 1333.700 ;
        RECT 1752.260 1331.900 1753.860 1333.700 ;
        RECT 1848.860 1331.900 1850.460 1333.700 ;
        RECT 1945.460 1331.900 1947.060 1333.700 ;
        RECT 2042.060 1331.900 2043.660 1333.700 ;
        RECT 2138.660 1331.900 2140.260 1333.700 ;
        RECT 2235.260 1331.900 2236.860 1333.700 ;
        RECT 2331.860 1331.900 2333.460 1333.700 ;
        RECT 2428.460 1331.900 2430.060 1333.700 ;
        RECT 2525.060 1331.900 2526.660 1333.700 ;
        RECT 2621.660 1331.900 2623.260 1337.100 ;
        RECT 1205.780 1330.300 1208.300 1331.900 ;
        RECT 1544.340 1330.300 1560.660 1331.900 ;
        RECT 1640.940 1330.300 1657.260 1331.900 ;
        RECT 1737.540 1330.300 1753.860 1331.900 ;
        RECT 1834.140 1330.300 1850.460 1331.900 ;
        RECT 1930.740 1330.300 1947.060 1331.900 ;
        RECT 2027.340 1330.300 2043.660 1331.900 ;
        RECT 2123.940 1330.300 2140.260 1331.900 ;
        RECT 2220.540 1330.300 2236.860 1331.900 ;
        RECT 2317.140 1330.300 2333.460 1331.900 ;
        RECT 2413.740 1330.300 2430.060 1331.900 ;
        RECT 2510.340 1330.300 2526.660 1331.900 ;
        RECT 2606.940 1330.300 2623.260 1331.900 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 943.070 1339.500 943.390 1339.560 ;
        RECT 2697.970 1339.500 2698.290 1339.560 ;
        RECT 943.070 1339.360 2698.290 1339.500 ;
        RECT 943.070 1339.300 943.390 1339.360 ;
        RECT 2697.970 1339.300 2698.290 1339.360 ;
      LAYER via ;
        RECT 943.100 1339.300 943.360 1339.560 ;
        RECT 2698.000 1339.300 2698.260 1339.560 ;
      LAYER met2 ;
        RECT 943.100 1339.270 943.360 1339.590 ;
        RECT 2698.000 1339.270 2698.260 1339.590 ;
        RECT 943.160 1325.025 943.300 1339.270 ;
        RECT 943.050 1321.025 943.330 1325.025 ;
        RECT 2698.060 17.410 2698.200 1339.270 ;
        RECT 2698.060 17.270 2702.800 17.410 ;
        RECT 2702.660 2.400 2702.800 17.270 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.010 1322.330 1047.290 1325.025 ;
        RECT 1048.430 1322.330 1048.710 1322.445 ;
        RECT 1047.010 1322.190 1048.710 1322.330 ;
        RECT 1047.010 1321.025 1047.290 1322.190 ;
        RECT 1048.430 1322.075 1048.710 1322.190 ;
        RECT 2718.690 1322.075 2718.970 1322.445 ;
        RECT 2718.760 17.410 2718.900 1322.075 ;
        RECT 2718.760 17.270 2720.740 17.410 ;
        RECT 2720.600 2.400 2720.740 17.270 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
      LAYER via2 ;
        RECT 1048.430 1322.120 1048.710 1322.400 ;
        RECT 2718.690 1322.120 2718.970 1322.400 ;
      LAYER met3 ;
        RECT 1048.405 1322.410 1048.735 1322.425 ;
        RECT 2718.665 1322.410 2718.995 1322.425 ;
        RECT 1048.405 1322.110 2718.995 1322.410 ;
        RECT 1048.405 1322.095 1048.735 1322.110 ;
        RECT 2718.665 1322.095 2718.995 1322.110 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.670 200.500 648.990 200.560 ;
        RECT 655.110 200.500 655.430 200.560 ;
        RECT 648.670 200.360 655.430 200.500 ;
        RECT 648.670 200.300 648.990 200.360 ;
        RECT 655.110 200.300 655.430 200.360 ;
        RECT 655.110 107.000 655.430 107.060 ;
        RECT 2732.930 107.000 2733.250 107.060 ;
        RECT 655.110 106.860 2733.250 107.000 ;
        RECT 655.110 106.800 655.430 106.860 ;
        RECT 2732.930 106.800 2733.250 106.860 ;
      LAYER via ;
        RECT 648.700 200.300 648.960 200.560 ;
        RECT 655.140 200.300 655.400 200.560 ;
        RECT 655.140 106.800 655.400 107.060 ;
        RECT 2732.960 106.800 2733.220 107.060 ;
      LAYER met2 ;
        RECT 648.650 216.000 648.930 220.000 ;
        RECT 648.760 200.590 648.900 216.000 ;
        RECT 648.700 200.270 648.960 200.590 ;
        RECT 655.140 200.270 655.400 200.590 ;
        RECT 655.200 107.090 655.340 200.270 ;
        RECT 655.140 106.770 655.400 107.090 ;
        RECT 2732.960 106.770 2733.220 107.090 ;
        RECT 2733.020 17.410 2733.160 106.770 ;
        RECT 2733.020 17.270 2738.680 17.410 ;
        RECT 2738.540 2.400 2738.680 17.270 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1393.410 25.060 1393.730 25.120 ;
        RECT 2755.930 25.060 2756.250 25.120 ;
        RECT 1393.410 24.920 2756.250 25.060 ;
        RECT 1393.410 24.860 1393.730 24.920 ;
        RECT 2755.930 24.860 2756.250 24.920 ;
      LAYER via ;
        RECT 1393.440 24.860 1393.700 25.120 ;
        RECT 2755.960 24.860 2756.220 25.120 ;
      LAYER met2 ;
        RECT 1390.170 216.650 1390.450 220.000 ;
        RECT 1390.170 216.510 1393.640 216.650 ;
        RECT 1390.170 216.000 1390.450 216.510 ;
        RECT 1393.500 25.150 1393.640 216.510 ;
        RECT 1393.440 24.830 1393.700 25.150 ;
        RECT 2755.960 24.830 2756.220 25.150 ;
        RECT 2756.020 2.400 2756.160 24.830 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 834.510 60.420 834.830 60.480 ;
        RECT 1235.170 60.420 1235.490 60.480 ;
        RECT 834.510 60.280 1235.490 60.420 ;
        RECT 834.510 60.220 834.830 60.280 ;
        RECT 1235.170 60.220 1235.490 60.280 ;
        RECT 829.450 14.860 829.770 14.920 ;
        RECT 834.510 14.860 834.830 14.920 ;
        RECT 829.450 14.720 834.830 14.860 ;
        RECT 829.450 14.660 829.770 14.720 ;
        RECT 834.510 14.660 834.830 14.720 ;
      LAYER via ;
        RECT 834.540 60.220 834.800 60.480 ;
        RECT 1235.200 60.220 1235.460 60.480 ;
        RECT 829.480 14.660 829.740 14.920 ;
        RECT 834.540 14.660 834.800 14.920 ;
      LAYER met2 ;
        RECT 1237.450 216.650 1237.730 220.000 ;
        RECT 1235.260 216.510 1237.730 216.650 ;
        RECT 1235.260 60.510 1235.400 216.510 ;
        RECT 1237.450 216.000 1237.730 216.510 ;
        RECT 834.540 60.190 834.800 60.510 ;
        RECT 1235.200 60.190 1235.460 60.510 ;
        RECT 834.600 14.950 834.740 60.190 ;
        RECT 829.480 14.630 829.740 14.950 ;
        RECT 834.540 14.630 834.800 14.950 ;
        RECT 829.540 2.400 829.680 14.630 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 1328.875 443.810 1329.245 ;
        RECT 2773.890 1328.875 2774.170 1329.245 ;
        RECT 443.600 1325.025 443.740 1328.875 ;
        RECT 443.490 1321.025 443.770 1325.025 ;
        RECT 2773.960 2.400 2774.100 1328.875 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
      LAYER via2 ;
        RECT 443.530 1328.920 443.810 1329.200 ;
        RECT 2773.890 1328.920 2774.170 1329.200 ;
      LAYER met3 ;
        RECT 443.505 1329.210 443.835 1329.225 ;
        RECT 2773.865 1329.210 2774.195 1329.225 ;
        RECT 443.505 1328.910 2774.195 1329.210 ;
        RECT 443.505 1328.895 443.835 1328.910 ;
        RECT 2773.865 1328.895 2774.195 1328.910 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2791.830 32.795 2792.110 33.165 ;
        RECT 2791.900 2.400 2792.040 32.795 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
      LAYER via2 ;
        RECT 2791.830 32.840 2792.110 33.120 ;
      LAYER met3 ;
        RECT 280.870 1061.290 281.250 1061.300 ;
        RECT 280.870 1061.200 310.500 1061.290 ;
        RECT 280.870 1060.990 314.000 1061.200 ;
        RECT 280.870 1060.980 281.250 1060.990 ;
        RECT 310.000 1060.600 314.000 1060.990 ;
        RECT 280.870 33.130 281.250 33.140 ;
        RECT 2791.805 33.130 2792.135 33.145 ;
        RECT 280.870 32.830 2792.135 33.130 ;
        RECT 280.870 32.820 281.250 32.830 ;
        RECT 2791.805 32.815 2792.135 32.830 ;
      LAYER via3 ;
        RECT 280.900 1060.980 281.220 1061.300 ;
        RECT 280.900 32.820 281.220 33.140 ;
      LAYER met4 ;
        RECT 280.895 1060.975 281.225 1061.305 ;
        RECT 280.910 33.145 281.210 1060.975 ;
        RECT 280.895 32.815 281.225 33.145 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 435.100 1419.490 435.160 ;
        RECT 1590.290 435.100 1590.610 435.160 ;
        RECT 1419.170 434.960 1590.610 435.100 ;
        RECT 1419.170 434.900 1419.490 434.960 ;
        RECT 1590.290 434.900 1590.610 434.960 ;
        RECT 1590.290 237.900 1590.610 237.960 ;
        RECT 2808.370 237.900 2808.690 237.960 ;
        RECT 1590.290 237.760 2808.690 237.900 ;
        RECT 1590.290 237.700 1590.610 237.760 ;
        RECT 2808.370 237.700 2808.690 237.760 ;
      LAYER via ;
        RECT 1419.200 434.900 1419.460 435.160 ;
        RECT 1590.320 434.900 1590.580 435.160 ;
        RECT 1590.320 237.700 1590.580 237.960 ;
        RECT 2808.400 237.700 2808.660 237.960 ;
      LAYER met2 ;
        RECT 1419.190 439.435 1419.470 439.805 ;
        RECT 1419.260 435.190 1419.400 439.435 ;
        RECT 1419.200 434.870 1419.460 435.190 ;
        RECT 1590.320 434.870 1590.580 435.190 ;
        RECT 1590.380 237.990 1590.520 434.870 ;
        RECT 1590.320 237.670 1590.580 237.990 ;
        RECT 2808.400 237.670 2808.660 237.990 ;
        RECT 2808.460 17.410 2808.600 237.670 ;
        RECT 2808.460 17.270 2809.980 17.410 ;
        RECT 2809.840 2.400 2809.980 17.270 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
      LAYER via2 ;
        RECT 1419.190 439.480 1419.470 439.760 ;
      LAYER met3 ;
        RECT 1419.165 439.770 1419.495 439.785 ;
        RECT 1408.060 439.680 1419.495 439.770 ;
        RECT 1404.305 439.470 1419.495 439.680 ;
        RECT 1404.305 439.080 1408.305 439.470 ;
        RECT 1419.165 439.455 1419.495 439.470 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2827.710 32.115 2827.990 32.485 ;
        RECT 2827.780 2.400 2827.920 32.115 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
      LAYER via2 ;
        RECT 2827.710 32.160 2827.990 32.440 ;
      LAYER met3 ;
        RECT 288.230 738.970 288.610 738.980 ;
        RECT 288.230 738.880 310.500 738.970 ;
        RECT 288.230 738.670 314.000 738.880 ;
        RECT 288.230 738.660 288.610 738.670 ;
        RECT 310.000 738.280 314.000 738.670 ;
        RECT 288.230 32.450 288.610 32.460 ;
        RECT 2827.685 32.450 2828.015 32.465 ;
        RECT 288.230 32.150 2828.015 32.450 ;
        RECT 288.230 32.140 288.610 32.150 ;
        RECT 2827.685 32.135 2828.015 32.150 ;
      LAYER via3 ;
        RECT 288.260 738.660 288.580 738.980 ;
        RECT 288.260 32.140 288.580 32.460 ;
      LAYER met4 ;
        RECT 288.255 738.655 288.585 738.985 ;
        RECT 288.270 32.465 288.570 738.655 ;
        RECT 288.255 32.135 288.585 32.465 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 280.210 586.740 280.530 586.800 ;
        RECT 296.770 586.740 297.090 586.800 ;
        RECT 280.210 586.600 297.090 586.740 ;
        RECT 280.210 586.540 280.530 586.600 ;
        RECT 296.770 586.540 297.090 586.600 ;
      LAYER via ;
        RECT 280.240 586.540 280.500 586.800 ;
        RECT 296.800 586.540 297.060 586.800 ;
      LAYER met2 ;
        RECT 296.790 593.115 297.070 593.485 ;
        RECT 296.860 586.830 297.000 593.115 ;
        RECT 280.240 586.510 280.500 586.830 ;
        RECT 296.800 586.510 297.060 586.830 ;
        RECT 280.300 31.805 280.440 586.510 ;
        RECT 280.230 31.435 280.510 31.805 ;
        RECT 2845.190 31.435 2845.470 31.805 ;
        RECT 2845.260 2.400 2845.400 31.435 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
      LAYER via2 ;
        RECT 296.790 593.160 297.070 593.440 ;
        RECT 280.230 31.480 280.510 31.760 ;
        RECT 2845.190 31.480 2845.470 31.760 ;
      LAYER met3 ;
        RECT 296.765 593.450 297.095 593.465 ;
        RECT 296.765 593.360 310.500 593.450 ;
        RECT 296.765 593.150 314.000 593.360 ;
        RECT 296.765 593.135 297.095 593.150 ;
        RECT 310.000 592.760 314.000 593.150 ;
        RECT 280.205 31.770 280.535 31.785 ;
        RECT 2845.165 31.770 2845.495 31.785 ;
        RECT 280.205 31.470 2845.495 31.770 ;
        RECT 280.205 31.455 280.535 31.470 ;
        RECT 2845.165 31.455 2845.495 31.470 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 286.190 648.960 286.510 649.020 ;
        RECT 298.610 648.960 298.930 649.020 ;
        RECT 286.190 648.820 298.930 648.960 ;
        RECT 286.190 648.760 286.510 648.820 ;
        RECT 298.610 648.760 298.930 648.820 ;
      LAYER via ;
        RECT 286.220 648.760 286.480 649.020 ;
        RECT 298.640 648.760 298.900 649.020 ;
      LAYER met2 ;
        RECT 298.630 651.595 298.910 651.965 ;
        RECT 298.700 649.050 298.840 651.595 ;
        RECT 286.220 648.730 286.480 649.050 ;
        RECT 298.640 648.730 298.900 649.050 ;
        RECT 286.280 31.125 286.420 648.730 ;
        RECT 286.210 30.755 286.490 31.125 ;
        RECT 2863.130 30.755 2863.410 31.125 ;
        RECT 2863.200 2.400 2863.340 30.755 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
      LAYER via2 ;
        RECT 298.630 651.640 298.910 651.920 ;
        RECT 286.210 30.800 286.490 31.080 ;
        RECT 2863.130 30.800 2863.410 31.080 ;
      LAYER met3 ;
        RECT 298.605 651.930 298.935 651.945 ;
        RECT 298.605 651.840 310.500 651.930 ;
        RECT 298.605 651.630 314.000 651.840 ;
        RECT 298.605 651.615 298.935 651.630 ;
        RECT 310.000 651.240 314.000 651.630 ;
        RECT 286.185 31.090 286.515 31.105 ;
        RECT 2863.105 31.090 2863.435 31.105 ;
        RECT 286.185 30.790 2863.435 31.090 ;
        RECT 286.185 30.775 286.515 30.790 ;
        RECT 2863.105 30.775 2863.435 30.790 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.250 1321.650 1274.530 1325.025 ;
        RECT 1275.670 1321.650 1275.950 1321.765 ;
        RECT 1274.250 1321.510 1275.950 1321.650 ;
        RECT 1274.250 1321.025 1274.530 1321.510 ;
        RECT 1275.670 1321.395 1275.950 1321.510 ;
        RECT 2877.390 1318.675 2877.670 1319.045 ;
        RECT 2877.460 17.410 2877.600 1318.675 ;
        RECT 2877.460 17.270 2881.280 17.410 ;
        RECT 2881.140 2.400 2881.280 17.270 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
      LAYER via2 ;
        RECT 1275.670 1321.440 1275.950 1321.720 ;
        RECT 2877.390 1318.720 2877.670 1319.000 ;
      LAYER met3 ;
        RECT 1275.645 1321.730 1275.975 1321.745 ;
        RECT 1295.630 1321.730 1296.010 1321.740 ;
        RECT 1275.645 1321.430 1296.010 1321.730 ;
        RECT 1275.645 1321.415 1275.975 1321.430 ;
        RECT 1295.630 1321.420 1296.010 1321.430 ;
        RECT 1295.630 1319.010 1296.010 1319.020 ;
        RECT 2877.365 1319.010 2877.695 1319.025 ;
        RECT 1295.630 1318.710 2877.695 1319.010 ;
        RECT 1295.630 1318.700 1296.010 1318.710 ;
        RECT 2877.365 1318.695 2877.695 1318.710 ;
      LAYER via3 ;
        RECT 1295.660 1321.420 1295.980 1321.740 ;
        RECT 1295.660 1318.700 1295.980 1319.020 ;
      LAYER met4 ;
        RECT 1295.655 1321.415 1295.985 1321.745 ;
        RECT 1295.670 1319.025 1295.970 1321.415 ;
        RECT 1295.655 1318.695 1295.985 1319.025 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 352.430 200.500 352.750 200.560 ;
        RECT 358.410 200.500 358.730 200.560 ;
        RECT 352.430 200.360 358.730 200.500 ;
        RECT 352.430 200.300 352.750 200.360 ;
        RECT 358.410 200.300 358.730 200.360 ;
        RECT 358.410 24.040 358.730 24.100 ;
        RECT 2898.990 24.040 2899.310 24.100 ;
        RECT 358.410 23.900 2899.310 24.040 ;
        RECT 358.410 23.840 358.730 23.900 ;
        RECT 2898.990 23.840 2899.310 23.900 ;
      LAYER via ;
        RECT 352.460 200.300 352.720 200.560 ;
        RECT 358.440 200.300 358.700 200.560 ;
        RECT 358.440 23.840 358.700 24.100 ;
        RECT 2899.020 23.840 2899.280 24.100 ;
      LAYER met2 ;
        RECT 352.410 216.000 352.690 220.000 ;
        RECT 352.520 200.590 352.660 216.000 ;
        RECT 352.460 200.270 352.720 200.590 ;
        RECT 358.440 200.270 358.700 200.590 ;
        RECT 358.500 24.130 358.640 200.270 ;
        RECT 358.440 23.810 358.700 24.130 ;
        RECT 2899.020 23.810 2899.280 24.130 ;
        RECT 2899.080 2.400 2899.220 23.810 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 817.030 200.500 817.350 200.560 ;
        RECT 820.710 200.500 821.030 200.560 ;
        RECT 817.030 200.360 821.030 200.500 ;
        RECT 817.030 200.300 817.350 200.360 ;
        RECT 820.710 200.300 821.030 200.360 ;
        RECT 820.710 165.820 821.030 165.880 ;
        RECT 841.870 165.820 842.190 165.880 ;
        RECT 820.710 165.680 842.190 165.820 ;
        RECT 820.710 165.620 821.030 165.680 ;
        RECT 841.870 165.620 842.190 165.680 ;
      LAYER via ;
        RECT 817.060 200.300 817.320 200.560 ;
        RECT 820.740 200.300 821.000 200.560 ;
        RECT 820.740 165.620 821.000 165.880 ;
        RECT 841.900 165.620 842.160 165.880 ;
      LAYER met2 ;
        RECT 817.010 216.000 817.290 220.000 ;
        RECT 817.120 200.590 817.260 216.000 ;
        RECT 817.060 200.270 817.320 200.590 ;
        RECT 820.740 200.270 821.000 200.590 ;
        RECT 820.800 165.910 820.940 200.270 ;
        RECT 820.740 165.590 821.000 165.910 ;
        RECT 841.900 165.590 842.160 165.910 ;
        RECT 841.960 17.410 842.100 165.590 ;
        RECT 841.960 17.270 847.160 17.410 ;
        RECT 847.020 2.400 847.160 17.270 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 1321.650 798.010 1321.765 ;
        RECT 799.530 1321.650 799.810 1325.025 ;
        RECT 797.730 1321.510 799.810 1321.650 ;
        RECT 797.730 1321.395 798.010 1321.510 ;
        RECT 799.530 1321.025 799.810 1321.510 ;
        RECT 864.890 34.155 865.170 34.525 ;
        RECT 864.960 2.400 865.100 34.155 ;
        RECT 864.750 -4.800 865.310 2.400 ;
      LAYER via2 ;
        RECT 797.730 1321.440 798.010 1321.720 ;
        RECT 864.890 34.200 865.170 34.480 ;
      LAYER met3 ;
        RECT 779.510 1321.730 779.890 1321.740 ;
        RECT 797.705 1321.730 798.035 1321.745 ;
        RECT 779.510 1321.430 798.035 1321.730 ;
        RECT 779.510 1321.420 779.890 1321.430 ;
        RECT 797.705 1321.415 798.035 1321.430 ;
        RECT 316.750 1318.330 317.130 1318.340 ;
        RECT 779.510 1318.330 779.890 1318.340 ;
        RECT 316.750 1318.030 779.890 1318.330 ;
        RECT 316.750 1318.020 317.130 1318.030 ;
        RECT 779.510 1318.020 779.890 1318.030 ;
        RECT 317.670 219.450 318.050 219.460 ;
        RECT 326.870 219.450 327.250 219.460 ;
        RECT 317.670 219.150 327.250 219.450 ;
        RECT 317.670 219.140 318.050 219.150 ;
        RECT 326.870 219.140 327.250 219.150 ;
        RECT 326.870 34.490 327.250 34.500 ;
        RECT 864.865 34.490 865.195 34.505 ;
        RECT 326.870 34.190 865.195 34.490 ;
        RECT 326.870 34.180 327.250 34.190 ;
        RECT 864.865 34.175 865.195 34.190 ;
      LAYER via3 ;
        RECT 779.540 1321.420 779.860 1321.740 ;
        RECT 316.780 1318.020 317.100 1318.340 ;
        RECT 779.540 1318.020 779.860 1318.340 ;
        RECT 317.700 219.140 318.020 219.460 ;
        RECT 326.900 219.140 327.220 219.460 ;
        RECT 326.900 34.180 327.220 34.500 ;
      LAYER met4 ;
        RECT 779.535 1321.415 779.865 1321.745 ;
        RECT 779.550 1318.345 779.850 1321.415 ;
        RECT 316.775 1318.015 317.105 1318.345 ;
        RECT 779.535 1318.015 779.865 1318.345 ;
        RECT 316.790 1201.370 317.090 1318.015 ;
        RECT 316.790 1201.070 318.010 1201.370 ;
        RECT 317.710 1198.650 318.010 1201.070 ;
        RECT 316.790 1198.350 318.010 1198.650 ;
        RECT 316.790 1195.250 317.090 1198.350 ;
        RECT 315.870 1194.950 317.090 1195.250 ;
        RECT 315.870 1110.250 316.170 1194.950 ;
        RECT 314.950 1109.950 316.170 1110.250 ;
        RECT 314.950 1103.450 315.250 1109.950 ;
        RECT 314.030 1103.150 315.250 1103.450 ;
        RECT 314.030 1061.290 314.330 1103.150 ;
        RECT 314.030 1060.990 318.010 1061.290 ;
        RECT 317.710 1055.850 318.010 1060.990 ;
        RECT 316.790 1055.550 318.010 1055.850 ;
        RECT 316.790 1008.250 317.090 1055.550 ;
        RECT 315.870 1007.950 317.090 1008.250 ;
        RECT 315.870 981.050 316.170 1007.950 ;
        RECT 315.870 980.750 318.010 981.050 ;
        RECT 317.710 953.850 318.010 980.750 ;
        RECT 317.710 953.550 321.690 953.850 ;
        RECT 321.390 916.450 321.690 953.550 ;
        RECT 320.470 916.150 321.690 916.450 ;
        RECT 320.470 913.050 320.770 916.150 ;
        RECT 319.550 912.750 320.770 913.050 ;
        RECT 319.550 885.850 319.850 912.750 ;
        RECT 316.790 885.550 319.850 885.850 ;
        RECT 316.790 868.850 317.090 885.550 ;
        RECT 316.790 868.550 318.010 868.850 ;
        RECT 317.710 770.250 318.010 868.550 ;
        RECT 315.870 769.950 318.010 770.250 ;
        RECT 315.870 746.450 316.170 769.950 ;
        RECT 315.870 746.150 318.010 746.450 ;
        RECT 317.710 641.050 318.010 746.150 ;
        RECT 316.790 640.750 318.010 641.050 ;
        RECT 316.790 627.450 317.090 640.750 ;
        RECT 316.790 627.150 318.930 627.450 ;
        RECT 318.630 579.850 318.930 627.150 ;
        RECT 316.790 579.550 318.930 579.850 ;
        RECT 316.790 552.650 317.090 579.550 ;
        RECT 314.950 552.350 317.090 552.650 ;
        RECT 314.950 511.850 315.250 552.350 ;
        RECT 314.950 511.550 316.170 511.850 ;
        RECT 315.870 505.050 316.170 511.550 ;
        RECT 315.870 504.750 318.010 505.050 ;
        RECT 317.710 484.650 318.010 504.750 ;
        RECT 315.870 484.350 318.010 484.650 ;
        RECT 315.870 469.010 316.170 484.350 ;
        RECT 315.870 468.710 318.930 469.010 ;
        RECT 318.630 437.050 318.930 468.710 ;
        RECT 316.790 436.750 318.930 437.050 ;
        RECT 316.790 420.050 317.090 436.750 ;
        RECT 316.790 419.750 318.010 420.050 ;
        RECT 317.710 352.050 318.010 419.750 ;
        RECT 316.790 351.750 318.010 352.050 ;
        RECT 316.790 243.250 317.090 351.750 ;
        RECT 316.790 242.950 318.010 243.250 ;
        RECT 317.710 219.465 318.010 242.950 ;
        RECT 317.695 219.135 318.025 219.465 ;
        RECT 326.895 219.135 327.225 219.465 ;
        RECT 326.910 34.505 327.210 219.135 ;
        RECT 326.895 34.175 327.225 34.505 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 427.945 1318.605 428.115 1321.495 ;
      LAYER mcon ;
        RECT 427.945 1321.325 428.115 1321.495 ;
      LAYER met1 ;
        RECT 427.870 1321.480 428.190 1321.540 ;
        RECT 427.675 1321.340 428.190 1321.480 ;
        RECT 427.870 1321.280 428.190 1321.340 ;
        RECT 282.050 1318.760 282.370 1318.820 ;
        RECT 427.885 1318.760 428.175 1318.805 ;
        RECT 282.050 1318.620 428.175 1318.760 ;
        RECT 282.050 1318.560 282.370 1318.620 ;
        RECT 427.885 1318.575 428.175 1318.620 ;
        RECT 282.050 19.960 282.370 20.020 ;
        RECT 882.350 19.960 882.670 20.020 ;
        RECT 282.050 19.820 882.670 19.960 ;
        RECT 282.050 19.760 282.370 19.820 ;
        RECT 882.350 19.760 882.670 19.820 ;
      LAYER via ;
        RECT 427.900 1321.280 428.160 1321.540 ;
        RECT 282.080 1318.560 282.340 1318.820 ;
        RECT 282.080 19.760 282.340 20.020 ;
        RECT 882.380 19.760 882.640 20.020 ;
      LAYER met2 ;
        RECT 428.770 1321.650 429.050 1325.025 ;
        RECT 427.960 1321.570 429.050 1321.650 ;
        RECT 427.900 1321.510 429.050 1321.570 ;
        RECT 427.900 1321.250 428.160 1321.510 ;
        RECT 428.770 1321.025 429.050 1321.510 ;
        RECT 282.080 1318.530 282.340 1318.850 ;
        RECT 282.140 20.050 282.280 1318.530 ;
        RECT 282.080 19.730 282.340 20.050 ;
        RECT 882.380 19.730 882.640 20.050 ;
        RECT 882.440 16.050 882.580 19.730 ;
        RECT 882.440 15.910 883.040 16.050 ;
        RECT 882.900 2.400 883.040 15.910 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 900.750 26.080 901.070 26.140 ;
        RECT 993.670 26.080 993.990 26.140 ;
        RECT 900.750 25.940 993.990 26.080 ;
        RECT 900.750 25.880 901.070 25.940 ;
        RECT 993.670 25.880 993.990 25.940 ;
      LAYER via ;
        RECT 900.780 25.880 901.040 26.140 ;
        RECT 993.700 25.880 993.960 26.140 ;
      LAYER met2 ;
        RECT 994.570 216.650 994.850 220.000 ;
        RECT 993.760 216.510 994.850 216.650 ;
        RECT 993.760 26.170 993.900 216.510 ;
        RECT 994.570 216.000 994.850 216.510 ;
        RECT 900.780 25.850 901.040 26.170 ;
        RECT 993.700 25.850 993.960 26.170 ;
        RECT 900.840 2.400 900.980 25.850 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1389.805 1321.325 1389.975 1323.195 ;
      LAYER mcon ;
        RECT 1389.805 1323.025 1389.975 1323.195 ;
      LAYER met1 ;
        RECT 1389.745 1323.180 1390.035 1323.225 ;
        RECT 1428.830 1323.180 1429.150 1323.240 ;
        RECT 1389.745 1323.040 1429.150 1323.180 ;
        RECT 1389.745 1322.995 1390.035 1323.040 ;
        RECT 1428.830 1322.980 1429.150 1323.040 ;
        RECT 1092.570 1321.280 1092.890 1321.540 ;
        RECT 1389.745 1321.480 1390.035 1321.525 ;
        RECT 1122.560 1321.340 1390.035 1321.480 ;
        RECT 1092.660 1321.140 1092.800 1321.280 ;
        RECT 1122.560 1321.140 1122.700 1321.340 ;
        RECT 1389.745 1321.295 1390.035 1321.340 ;
        RECT 1092.660 1321.000 1122.700 1321.140 ;
        RECT 918.690 19.960 919.010 20.020 ;
        RECT 1428.830 19.960 1429.150 20.020 ;
        RECT 918.690 19.820 1429.150 19.960 ;
        RECT 918.690 19.760 919.010 19.820 ;
        RECT 1428.830 19.760 1429.150 19.820 ;
      LAYER via ;
        RECT 1428.860 1322.980 1429.120 1323.240 ;
        RECT 1092.600 1321.280 1092.860 1321.540 ;
        RECT 918.720 19.760 918.980 20.020 ;
        RECT 1428.860 19.760 1429.120 20.020 ;
      LAYER met2 ;
        RECT 1091.170 1321.650 1091.450 1325.025 ;
        RECT 1428.860 1322.950 1429.120 1323.270 ;
        RECT 1091.170 1321.570 1092.800 1321.650 ;
        RECT 1091.170 1321.510 1092.860 1321.570 ;
        RECT 1091.170 1321.025 1091.450 1321.510 ;
        RECT 1092.600 1321.250 1092.860 1321.510 ;
        RECT 1428.920 20.050 1429.060 1322.950 ;
        RECT 918.720 19.730 918.980 20.050 ;
        RECT 1428.860 19.730 1429.120 20.050 ;
        RECT 918.780 2.400 918.920 19.730 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.590 197.100 304.910 197.160 ;
        RECT 931.570 197.100 931.890 197.160 ;
        RECT 304.590 196.960 931.890 197.100 ;
        RECT 304.590 196.900 304.910 196.960 ;
        RECT 931.570 196.900 931.890 196.960 ;
        RECT 931.570 2.960 931.890 3.020 ;
        RECT 936.170 2.960 936.490 3.020 ;
        RECT 931.570 2.820 936.490 2.960 ;
        RECT 931.570 2.760 931.890 2.820 ;
        RECT 936.170 2.760 936.490 2.820 ;
      LAYER via ;
        RECT 304.620 196.900 304.880 197.160 ;
        RECT 931.600 196.900 931.860 197.160 ;
        RECT 931.600 2.760 931.860 3.020 ;
        RECT 936.200 2.760 936.460 3.020 ;
      LAYER met2 ;
        RECT 304.610 1097.675 304.890 1098.045 ;
        RECT 304.680 197.190 304.820 1097.675 ;
        RECT 304.620 196.870 304.880 197.190 ;
        RECT 931.600 196.870 931.860 197.190 ;
        RECT 931.660 3.050 931.800 196.870 ;
        RECT 931.600 2.730 931.860 3.050 ;
        RECT 936.200 2.730 936.460 3.050 ;
        RECT 936.260 2.400 936.400 2.730 ;
        RECT 936.050 -4.800 936.610 2.400 ;
      LAYER via2 ;
        RECT 304.610 1097.720 304.890 1098.000 ;
      LAYER met3 ;
        RECT 304.585 1098.010 304.915 1098.025 ;
        RECT 304.585 1097.920 310.500 1098.010 ;
        RECT 304.585 1097.710 314.000 1097.920 ;
        RECT 304.585 1097.695 304.915 1097.710 ;
        RECT 310.000 1097.320 314.000 1097.710 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 285.730 559.200 286.050 559.260 ;
        RECT 298.150 559.200 298.470 559.260 ;
        RECT 285.730 559.060 298.470 559.200 ;
        RECT 285.730 559.000 286.050 559.060 ;
        RECT 298.150 559.000 298.470 559.060 ;
        RECT 285.730 19.280 286.050 19.340 ;
        RECT 954.110 19.280 954.430 19.340 ;
        RECT 285.730 19.140 954.430 19.280 ;
        RECT 285.730 19.080 286.050 19.140 ;
        RECT 954.110 19.080 954.430 19.140 ;
      LAYER via ;
        RECT 285.760 559.000 286.020 559.260 ;
        RECT 298.180 559.000 298.440 559.260 ;
        RECT 285.760 19.080 286.020 19.340 ;
        RECT 954.140 19.080 954.400 19.340 ;
      LAYER met2 ;
        RECT 298.170 563.195 298.450 563.565 ;
        RECT 298.240 559.290 298.380 563.195 ;
        RECT 285.760 558.970 286.020 559.290 ;
        RECT 298.180 558.970 298.440 559.290 ;
        RECT 285.820 19.370 285.960 558.970 ;
        RECT 285.760 19.050 286.020 19.370 ;
        RECT 954.140 19.050 954.400 19.370 ;
        RECT 954.200 2.400 954.340 19.050 ;
        RECT 953.990 -4.800 954.550 2.400 ;
      LAYER via2 ;
        RECT 298.170 563.240 298.450 563.520 ;
      LAYER met3 ;
        RECT 298.145 563.530 298.475 563.545 ;
        RECT 298.145 563.440 310.500 563.530 ;
        RECT 298.145 563.230 314.000 563.440 ;
        RECT 298.145 563.215 298.475 563.230 ;
        RECT 310.000 562.840 314.000 563.230 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 306.890 189.960 307.210 190.020 ;
        RECT 966.070 189.960 966.390 190.020 ;
        RECT 306.890 189.820 966.390 189.960 ;
        RECT 306.890 189.760 307.210 189.820 ;
        RECT 966.070 189.760 966.390 189.820 ;
        RECT 966.070 14.520 966.390 14.580 ;
        RECT 972.050 14.520 972.370 14.580 ;
        RECT 966.070 14.380 972.370 14.520 ;
        RECT 966.070 14.320 966.390 14.380 ;
        RECT 972.050 14.320 972.370 14.380 ;
      LAYER via ;
        RECT 306.920 189.760 307.180 190.020 ;
        RECT 966.100 189.760 966.360 190.020 ;
        RECT 966.100 14.320 966.360 14.580 ;
        RECT 972.080 14.320 972.340 14.580 ;
      LAYER met2 ;
        RECT 306.910 431.275 307.190 431.645 ;
        RECT 306.980 190.050 307.120 431.275 ;
        RECT 306.920 189.730 307.180 190.050 ;
        RECT 966.100 189.730 966.360 190.050 ;
        RECT 966.160 14.610 966.300 189.730 ;
        RECT 966.100 14.290 966.360 14.610 ;
        RECT 972.080 14.290 972.340 14.610 ;
        RECT 972.140 2.400 972.280 14.290 ;
        RECT 971.930 -4.800 972.490 2.400 ;
      LAYER via2 ;
        RECT 306.910 431.320 307.190 431.600 ;
      LAYER met3 ;
        RECT 306.885 431.610 307.215 431.625 ;
        RECT 306.885 431.520 310.500 431.610 ;
        RECT 306.885 431.310 314.000 431.520 ;
        RECT 306.885 431.295 307.215 431.310 ;
        RECT 310.000 430.920 314.000 431.310 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 407.245 1318.945 407.415 1321.495 ;
        RECT 544.785 16.405 545.415 16.575 ;
      LAYER mcon ;
        RECT 407.245 1321.325 407.415 1321.495 ;
        RECT 545.245 16.405 545.415 16.575 ;
      LAYER met1 ;
        RECT 407.170 1321.480 407.490 1321.540 ;
        RECT 406.975 1321.340 407.490 1321.480 ;
        RECT 407.170 1321.280 407.490 1321.340 ;
        RECT 282.510 1319.100 282.830 1319.160 ;
        RECT 407.185 1319.100 407.475 1319.145 ;
        RECT 282.510 1318.960 407.475 1319.100 ;
        RECT 282.510 1318.900 282.830 1318.960 ;
        RECT 407.185 1318.915 407.475 1318.960 ;
        RECT 282.510 16.560 282.830 16.620 ;
        RECT 544.725 16.560 545.015 16.605 ;
        RECT 282.510 16.420 545.015 16.560 ;
        RECT 282.510 16.360 282.830 16.420 ;
        RECT 544.725 16.375 545.015 16.420 ;
        RECT 545.185 16.560 545.475 16.605 ;
        RECT 545.185 16.420 632.800 16.560 ;
        RECT 545.185 16.375 545.475 16.420 ;
        RECT 632.660 15.880 632.800 16.420 ;
        RECT 650.970 15.880 651.290 15.940 ;
        RECT 632.660 15.740 651.290 15.880 ;
        RECT 650.970 15.680 651.290 15.740 ;
      LAYER via ;
        RECT 407.200 1321.280 407.460 1321.540 ;
        RECT 282.540 1318.900 282.800 1319.160 ;
        RECT 282.540 16.360 282.800 16.620 ;
        RECT 651.000 15.680 651.260 15.940 ;
      LAYER met2 ;
        RECT 408.530 1321.650 408.810 1325.025 ;
        RECT 407.260 1321.570 408.810 1321.650 ;
        RECT 407.200 1321.510 408.810 1321.570 ;
        RECT 407.200 1321.250 407.460 1321.510 ;
        RECT 408.530 1321.025 408.810 1321.510 ;
        RECT 282.540 1318.870 282.800 1319.190 ;
        RECT 282.600 16.650 282.740 1318.870 ;
        RECT 282.540 16.330 282.800 16.650 ;
        RECT 651.000 15.650 651.260 15.970 ;
        RECT 651.060 2.400 651.200 15.650 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 288.490 1335.080 288.810 1335.140 ;
        RECT 581.510 1335.080 581.830 1335.140 ;
        RECT 288.490 1334.940 581.830 1335.080 ;
        RECT 288.490 1334.880 288.810 1334.940 ;
        RECT 581.510 1334.880 581.830 1334.940 ;
        RECT 288.490 18.260 288.810 18.320 ;
        RECT 989.990 18.260 990.310 18.320 ;
        RECT 288.490 18.120 990.310 18.260 ;
        RECT 288.490 18.060 288.810 18.120 ;
        RECT 989.990 18.060 990.310 18.120 ;
      LAYER via ;
        RECT 288.520 1334.880 288.780 1335.140 ;
        RECT 581.540 1334.880 581.800 1335.140 ;
        RECT 288.520 18.060 288.780 18.320 ;
        RECT 990.020 18.060 990.280 18.320 ;
      LAYER met2 ;
        RECT 288.520 1334.850 288.780 1335.170 ;
        RECT 581.540 1334.850 581.800 1335.170 ;
        RECT 288.580 18.350 288.720 1334.850 ;
        RECT 581.600 1325.025 581.740 1334.850 ;
        RECT 581.490 1321.025 581.770 1325.025 ;
        RECT 288.520 18.030 288.780 18.350 ;
        RECT 990.020 18.030 990.280 18.350 ;
        RECT 990.080 2.400 990.220 18.030 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 662.010 25.400 662.330 25.460 ;
        RECT 1007.470 25.400 1007.790 25.460 ;
        RECT 662.010 25.260 1007.790 25.400 ;
        RECT 662.010 25.200 662.330 25.260 ;
        RECT 1007.470 25.200 1007.790 25.260 ;
      LAYER via ;
        RECT 662.040 25.200 662.300 25.460 ;
        RECT 1007.500 25.200 1007.760 25.460 ;
      LAYER met2 ;
        RECT 658.770 216.650 659.050 220.000 ;
        RECT 658.770 216.510 662.240 216.650 ;
        RECT 658.770 216.000 659.050 216.510 ;
        RECT 662.100 25.490 662.240 216.510 ;
        RECT 662.040 25.170 662.300 25.490 ;
        RECT 1007.500 25.170 1007.760 25.490 ;
        RECT 1007.560 2.400 1007.700 25.170 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1390.265 1322.005 1390.435 1322.855 ;
      LAYER mcon ;
        RECT 1390.265 1322.685 1390.435 1322.855 ;
      LAYER met1 ;
        RECT 1390.205 1322.840 1390.495 1322.885 ;
        RECT 1423.310 1322.840 1423.630 1322.900 ;
        RECT 1390.205 1322.700 1423.630 1322.840 ;
        RECT 1390.205 1322.655 1390.495 1322.700 ;
        RECT 1423.310 1322.640 1423.630 1322.700 ;
        RECT 1041.970 1322.160 1042.290 1322.220 ;
        RECT 1390.205 1322.160 1390.495 1322.205 ;
        RECT 1041.970 1322.020 1390.495 1322.160 ;
        RECT 1041.970 1321.960 1042.290 1322.020 ;
        RECT 1390.205 1321.975 1390.495 1322.020 ;
        RECT 1397.090 207.300 1397.410 207.360 ;
        RECT 1423.310 207.300 1423.630 207.360 ;
        RECT 1397.090 207.160 1423.630 207.300 ;
        RECT 1397.090 207.100 1397.410 207.160 ;
        RECT 1423.310 207.100 1423.630 207.160 ;
        RECT 1025.410 20.300 1025.730 20.360 ;
        RECT 1397.090 20.300 1397.410 20.360 ;
        RECT 1025.410 20.160 1397.410 20.300 ;
        RECT 1025.410 20.100 1025.730 20.160 ;
        RECT 1397.090 20.100 1397.410 20.160 ;
      LAYER via ;
        RECT 1423.340 1322.640 1423.600 1322.900 ;
        RECT 1042.000 1321.960 1042.260 1322.220 ;
        RECT 1397.120 207.100 1397.380 207.360 ;
        RECT 1423.340 207.100 1423.600 207.360 ;
        RECT 1025.440 20.100 1025.700 20.360 ;
        RECT 1397.120 20.100 1397.380 20.360 ;
      LAYER met2 ;
        RECT 1041.490 1322.330 1041.770 1325.025 ;
        RECT 1423.340 1322.610 1423.600 1322.930 ;
        RECT 1041.490 1322.250 1042.200 1322.330 ;
        RECT 1041.490 1322.190 1042.260 1322.250 ;
        RECT 1041.490 1321.025 1041.770 1322.190 ;
        RECT 1042.000 1321.930 1042.260 1322.190 ;
        RECT 1423.400 207.390 1423.540 1322.610 ;
        RECT 1397.120 207.070 1397.380 207.390 ;
        RECT 1423.340 207.070 1423.600 207.390 ;
        RECT 1397.180 20.390 1397.320 207.070 ;
        RECT 1025.440 20.070 1025.700 20.390 ;
        RECT 1397.120 20.070 1397.380 20.390 ;
        RECT 1025.500 2.400 1025.640 20.070 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1043.350 25.400 1043.670 25.460 ;
        RECT 1304.170 25.400 1304.490 25.460 ;
        RECT 1043.350 25.260 1304.490 25.400 ;
        RECT 1043.350 25.200 1043.670 25.260 ;
        RECT 1304.170 25.200 1304.490 25.260 ;
      LAYER via ;
        RECT 1043.380 25.200 1043.640 25.460 ;
        RECT 1304.200 25.200 1304.460 25.460 ;
      LAYER met2 ;
        RECT 1306.450 216.650 1306.730 220.000 ;
        RECT 1304.260 216.510 1306.730 216.650 ;
        RECT 1304.260 25.490 1304.400 216.510 ;
        RECT 1306.450 216.000 1306.730 216.510 ;
        RECT 1043.380 25.170 1043.640 25.490 ;
        RECT 1304.200 25.170 1304.460 25.490 ;
        RECT 1043.440 2.400 1043.580 25.170 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 749.870 1326.920 750.190 1326.980 ;
        RECT 1422.850 1326.920 1423.170 1326.980 ;
        RECT 749.870 1326.780 1423.170 1326.920 ;
        RECT 749.870 1326.720 750.190 1326.780 ;
        RECT 1422.850 1326.720 1423.170 1326.780 ;
        RECT 1061.290 34.240 1061.610 34.300 ;
        RECT 1422.850 34.240 1423.170 34.300 ;
        RECT 1061.290 34.100 1423.170 34.240 ;
        RECT 1061.290 34.040 1061.610 34.100 ;
        RECT 1422.850 34.040 1423.170 34.100 ;
      LAYER via ;
        RECT 749.900 1326.720 750.160 1326.980 ;
        RECT 1422.880 1326.720 1423.140 1326.980 ;
        RECT 1061.320 34.040 1061.580 34.300 ;
        RECT 1422.880 34.040 1423.140 34.300 ;
      LAYER met2 ;
        RECT 749.900 1326.690 750.160 1327.010 ;
        RECT 1422.880 1326.690 1423.140 1327.010 ;
        RECT 749.960 1325.025 750.100 1326.690 ;
        RECT 749.850 1321.025 750.130 1325.025 ;
        RECT 1422.940 34.330 1423.080 1326.690 ;
        RECT 1061.320 34.010 1061.580 34.330 ;
        RECT 1422.880 34.010 1423.140 34.330 ;
        RECT 1061.380 2.400 1061.520 34.010 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 917.310 25.740 917.630 25.800 ;
        RECT 1079.230 25.740 1079.550 25.800 ;
        RECT 917.310 25.600 1079.550 25.740 ;
        RECT 917.310 25.540 917.630 25.600 ;
        RECT 1079.230 25.540 1079.550 25.600 ;
      LAYER via ;
        RECT 917.340 25.540 917.600 25.800 ;
        RECT 1079.260 25.540 1079.520 25.800 ;
      LAYER met2 ;
        RECT 915.450 216.650 915.730 220.000 ;
        RECT 915.450 216.510 917.540 216.650 ;
        RECT 915.450 216.000 915.730 216.510 ;
        RECT 917.400 25.830 917.540 216.510 ;
        RECT 917.340 25.510 917.600 25.830 ;
        RECT 1079.260 25.510 1079.520 25.830 ;
        RECT 1079.320 2.400 1079.460 25.510 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1096.710 169.560 1097.030 169.620 ;
        RECT 1411.810 169.560 1412.130 169.620 ;
        RECT 1096.710 169.420 1412.130 169.560 ;
        RECT 1096.710 169.360 1097.030 169.420 ;
        RECT 1411.810 169.360 1412.130 169.420 ;
      LAYER via ;
        RECT 1096.740 169.360 1097.000 169.620 ;
        RECT 1411.840 169.360 1412.100 169.620 ;
      LAYER met2 ;
        RECT 1411.830 461.195 1412.110 461.565 ;
        RECT 1411.900 169.650 1412.040 461.195 ;
        RECT 1096.740 169.330 1097.000 169.650 ;
        RECT 1411.840 169.330 1412.100 169.650 ;
        RECT 1096.800 2.400 1096.940 169.330 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
      LAYER via2 ;
        RECT 1411.830 461.240 1412.110 461.520 ;
      LAYER met3 ;
        RECT 1411.805 461.530 1412.135 461.545 ;
        RECT 1408.060 461.440 1412.135 461.530 ;
        RECT 1404.305 461.230 1412.135 461.440 ;
        RECT 1404.305 460.840 1408.305 461.230 ;
        RECT 1411.805 461.215 1412.135 461.230 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 288.030 911.100 288.350 911.160 ;
        RECT 299.530 911.100 299.850 911.160 ;
        RECT 288.030 910.960 299.850 911.100 ;
        RECT 288.030 910.900 288.350 910.960 ;
        RECT 299.530 910.900 299.850 910.960 ;
        RECT 288.030 18.940 288.350 19.000 ;
        RECT 1114.650 18.940 1114.970 19.000 ;
        RECT 288.030 18.800 1114.970 18.940 ;
        RECT 288.030 18.740 288.350 18.800 ;
        RECT 1114.650 18.740 1114.970 18.800 ;
      LAYER via ;
        RECT 288.060 910.900 288.320 911.160 ;
        RECT 299.560 910.900 299.820 911.160 ;
        RECT 288.060 18.740 288.320 19.000 ;
        RECT 1114.680 18.740 1114.940 19.000 ;
      LAYER met2 ;
        RECT 299.550 914.075 299.830 914.445 ;
        RECT 299.620 911.190 299.760 914.075 ;
        RECT 288.060 910.870 288.320 911.190 ;
        RECT 299.560 910.870 299.820 911.190 ;
        RECT 288.120 19.030 288.260 910.870 ;
        RECT 288.060 18.710 288.320 19.030 ;
        RECT 1114.680 18.710 1114.940 19.030 ;
        RECT 1114.740 2.400 1114.880 18.710 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
      LAYER via2 ;
        RECT 299.550 914.120 299.830 914.400 ;
      LAYER met3 ;
        RECT 299.525 914.410 299.855 914.425 ;
        RECT 299.525 914.320 310.500 914.410 ;
        RECT 299.525 914.110 314.000 914.320 ;
        RECT 299.525 914.095 299.855 914.110 ;
        RECT 310.000 913.720 314.000 914.110 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 731.010 155.620 731.330 155.680 ;
        RECT 1131.670 155.620 1131.990 155.680 ;
        RECT 731.010 155.480 1131.990 155.620 ;
        RECT 731.010 155.420 731.330 155.480 ;
        RECT 1131.670 155.420 1131.990 155.480 ;
      LAYER via ;
        RECT 731.040 155.420 731.300 155.680 ;
        RECT 1131.700 155.420 1131.960 155.680 ;
      LAYER met2 ;
        RECT 727.770 216.650 728.050 220.000 ;
        RECT 727.770 216.510 731.240 216.650 ;
        RECT 727.770 216.000 728.050 216.510 ;
        RECT 731.100 155.710 731.240 216.510 ;
        RECT 731.040 155.390 731.300 155.710 ;
        RECT 1131.700 155.390 1131.960 155.710 ;
        RECT 1131.760 17.410 1131.900 155.390 ;
        RECT 1131.760 17.270 1132.820 17.410 ;
        RECT 1132.680 2.400 1132.820 17.270 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1104.070 200.500 1104.390 200.560 ;
        RECT 1110.510 200.500 1110.830 200.560 ;
        RECT 1104.070 200.360 1110.830 200.500 ;
        RECT 1104.070 200.300 1104.390 200.360 ;
        RECT 1110.510 200.300 1110.830 200.360 ;
        RECT 1110.510 25.740 1110.830 25.800 ;
        RECT 1150.530 25.740 1150.850 25.800 ;
        RECT 1110.510 25.600 1150.850 25.740 ;
        RECT 1110.510 25.540 1110.830 25.600 ;
        RECT 1150.530 25.540 1150.850 25.600 ;
      LAYER via ;
        RECT 1104.100 200.300 1104.360 200.560 ;
        RECT 1110.540 200.300 1110.800 200.560 ;
        RECT 1110.540 25.540 1110.800 25.800 ;
        RECT 1150.560 25.540 1150.820 25.800 ;
      LAYER met2 ;
        RECT 1104.050 216.000 1104.330 220.000 ;
        RECT 1104.160 200.590 1104.300 216.000 ;
        RECT 1104.100 200.270 1104.360 200.590 ;
        RECT 1110.540 200.270 1110.800 200.590 ;
        RECT 1110.600 25.830 1110.740 200.270 ;
        RECT 1110.540 25.510 1110.800 25.830 ;
        RECT 1150.560 25.510 1150.820 25.830 ;
        RECT 1150.620 2.400 1150.760 25.510 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1188.250 159.160 1188.570 159.420 ;
        RECT 1188.340 158.740 1188.480 159.160 ;
        RECT 1188.250 158.480 1188.570 158.740 ;
        RECT 1187.330 62.460 1187.650 62.520 ;
        RECT 1188.710 62.460 1189.030 62.520 ;
        RECT 1187.330 62.320 1189.030 62.460 ;
        RECT 1187.330 62.260 1187.650 62.320 ;
        RECT 1188.710 62.260 1189.030 62.320 ;
        RECT 667.990 59.400 668.310 59.460 ;
        RECT 1187.330 59.400 1187.650 59.460 ;
        RECT 667.990 59.260 1187.650 59.400 ;
        RECT 667.990 59.200 668.310 59.260 ;
        RECT 1187.330 59.200 1187.650 59.260 ;
      LAYER via ;
        RECT 1188.280 159.160 1188.540 159.420 ;
        RECT 1188.280 158.480 1188.540 158.740 ;
        RECT 1187.360 62.260 1187.620 62.520 ;
        RECT 1188.740 62.260 1189.000 62.520 ;
        RECT 668.020 59.200 668.280 59.460 ;
        RECT 1187.360 59.200 1187.620 59.460 ;
      LAYER met2 ;
        RECT 1192.370 217.330 1192.650 220.000 ;
        RECT 1188.340 217.190 1192.650 217.330 ;
        RECT 1188.340 159.450 1188.480 217.190 ;
        RECT 1192.370 216.000 1192.650 217.190 ;
        RECT 1188.280 159.130 1188.540 159.450 ;
        RECT 1188.280 158.450 1188.540 158.770 ;
        RECT 1188.340 110.570 1188.480 158.450 ;
        RECT 1188.340 110.430 1188.940 110.570 ;
        RECT 1188.800 62.550 1188.940 110.430 ;
        RECT 1187.360 62.230 1187.620 62.550 ;
        RECT 1188.740 62.230 1189.000 62.550 ;
        RECT 1187.420 59.490 1187.560 62.230 ;
        RECT 668.020 59.170 668.280 59.490 ;
        RECT 1187.360 59.170 1187.620 59.490 ;
        RECT 668.080 14.010 668.220 59.170 ;
        RECT 668.080 13.870 669.140 14.010 ;
        RECT 669.000 2.400 669.140 13.870 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 421.430 200.500 421.750 200.560 ;
        RECT 427.410 200.500 427.730 200.560 ;
        RECT 421.430 200.360 427.730 200.500 ;
        RECT 421.430 200.300 421.750 200.360 ;
        RECT 427.410 200.300 427.730 200.360 ;
        RECT 427.410 121.960 427.730 122.020 ;
        RECT 1166.170 121.960 1166.490 122.020 ;
        RECT 427.410 121.820 1166.490 121.960 ;
        RECT 427.410 121.760 427.730 121.820 ;
        RECT 1166.170 121.760 1166.490 121.820 ;
      LAYER via ;
        RECT 421.460 200.300 421.720 200.560 ;
        RECT 427.440 200.300 427.700 200.560 ;
        RECT 427.440 121.760 427.700 122.020 ;
        RECT 1166.200 121.760 1166.460 122.020 ;
      LAYER met2 ;
        RECT 421.410 216.000 421.690 220.000 ;
        RECT 421.520 200.590 421.660 216.000 ;
        RECT 421.460 200.270 421.720 200.590 ;
        RECT 427.440 200.270 427.700 200.590 ;
        RECT 427.500 122.050 427.640 200.270 ;
        RECT 427.440 121.730 427.700 122.050 ;
        RECT 1166.200 121.730 1166.460 122.050 ;
        RECT 1166.260 17.410 1166.400 121.730 ;
        RECT 1166.260 17.270 1168.700 17.410 ;
        RECT 1168.560 2.400 1168.700 17.270 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 357.950 73.000 358.270 73.060 ;
        RECT 1180.430 73.000 1180.750 73.060 ;
        RECT 357.950 72.860 1180.750 73.000 ;
        RECT 357.950 72.800 358.270 72.860 ;
        RECT 1180.430 72.800 1180.750 72.860 ;
        RECT 1180.430 2.960 1180.750 3.020 ;
        RECT 1185.950 2.960 1186.270 3.020 ;
        RECT 1180.430 2.820 1186.270 2.960 ;
        RECT 1180.430 2.760 1180.750 2.820 ;
        RECT 1185.950 2.760 1186.270 2.820 ;
      LAYER via ;
        RECT 357.980 72.800 358.240 73.060 ;
        RECT 1180.460 72.800 1180.720 73.060 ;
        RECT 1180.460 2.760 1180.720 3.020 ;
        RECT 1185.980 2.760 1186.240 3.020 ;
      LAYER met2 ;
        RECT 357.010 216.650 357.290 220.000 ;
        RECT 357.010 216.510 358.180 216.650 ;
        RECT 357.010 216.000 357.290 216.510 ;
        RECT 358.040 73.090 358.180 216.510 ;
        RECT 357.980 72.770 358.240 73.090 ;
        RECT 1180.460 72.770 1180.720 73.090 ;
        RECT 1180.520 3.050 1180.660 72.770 ;
        RECT 1180.460 2.730 1180.720 3.050 ;
        RECT 1185.980 2.730 1186.240 3.050 ;
        RECT 1186.040 2.400 1186.180 2.730 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1407.670 190.640 1407.990 190.700 ;
        RECT 1392.580 190.500 1407.990 190.640 ;
        RECT 1207.110 190.300 1207.430 190.360 ;
        RECT 1392.580 190.300 1392.720 190.500 ;
        RECT 1407.670 190.440 1407.990 190.500 ;
        RECT 1207.110 190.160 1392.720 190.300 ;
        RECT 1207.110 190.100 1207.430 190.160 ;
        RECT 1203.890 16.560 1204.210 16.620 ;
        RECT 1207.110 16.560 1207.430 16.620 ;
        RECT 1203.890 16.420 1207.430 16.560 ;
        RECT 1203.890 16.360 1204.210 16.420 ;
        RECT 1207.110 16.360 1207.430 16.420 ;
      LAYER via ;
        RECT 1207.140 190.100 1207.400 190.360 ;
        RECT 1407.700 190.440 1407.960 190.700 ;
        RECT 1203.920 16.360 1204.180 16.620 ;
        RECT 1207.140 16.360 1207.400 16.620 ;
      LAYER met2 ;
        RECT 1407.690 326.555 1407.970 326.925 ;
        RECT 1407.760 190.730 1407.900 326.555 ;
        RECT 1407.700 190.410 1407.960 190.730 ;
        RECT 1207.140 190.070 1207.400 190.390 ;
        RECT 1207.200 16.650 1207.340 190.070 ;
        RECT 1203.920 16.330 1204.180 16.650 ;
        RECT 1207.140 16.330 1207.400 16.650 ;
        RECT 1203.980 2.400 1204.120 16.330 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
      LAYER via2 ;
        RECT 1407.690 326.600 1407.970 326.880 ;
      LAYER met3 ;
        RECT 1404.305 328.920 1408.305 329.520 ;
        RECT 1407.910 326.905 1408.210 328.920 ;
        RECT 1407.665 326.590 1408.210 326.905 ;
        RECT 1407.665 326.575 1407.995 326.590 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 267.790 1104.220 268.110 1104.280 ;
        RECT 296.770 1104.220 297.090 1104.280 ;
        RECT 267.790 1104.080 297.090 1104.220 ;
        RECT 267.790 1104.020 268.110 1104.080 ;
        RECT 296.770 1104.020 297.090 1104.080 ;
        RECT 267.790 18.600 268.110 18.660 ;
        RECT 1221.830 18.600 1222.150 18.660 ;
        RECT 267.790 18.460 1222.150 18.600 ;
        RECT 267.790 18.400 268.110 18.460 ;
        RECT 1221.830 18.400 1222.150 18.460 ;
      LAYER via ;
        RECT 267.820 1104.020 268.080 1104.280 ;
        RECT 296.800 1104.020 297.060 1104.280 ;
        RECT 267.820 18.400 268.080 18.660 ;
        RECT 1221.860 18.400 1222.120 18.660 ;
      LAYER met2 ;
        RECT 296.790 1104.475 297.070 1104.845 ;
        RECT 296.860 1104.310 297.000 1104.475 ;
        RECT 267.820 1103.990 268.080 1104.310 ;
        RECT 296.800 1103.990 297.060 1104.310 ;
        RECT 267.880 18.690 268.020 1103.990 ;
        RECT 267.820 18.370 268.080 18.690 ;
        RECT 1221.860 18.370 1222.120 18.690 ;
        RECT 1221.920 2.400 1222.060 18.370 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
      LAYER via2 ;
        RECT 296.790 1104.520 297.070 1104.800 ;
      LAYER met3 ;
        RECT 296.765 1104.810 297.095 1104.825 ;
        RECT 296.765 1104.720 310.500 1104.810 ;
        RECT 296.765 1104.510 314.000 1104.720 ;
        RECT 296.765 1104.495 297.095 1104.510 ;
        RECT 310.000 1104.120 314.000 1104.510 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.010 80.480 593.330 80.540 ;
        RECT 1235.630 80.480 1235.950 80.540 ;
        RECT 593.010 80.340 1235.950 80.480 ;
        RECT 593.010 80.280 593.330 80.340 ;
        RECT 1235.630 80.280 1235.950 80.340 ;
      LAYER via ;
        RECT 593.040 80.280 593.300 80.540 ;
        RECT 1235.660 80.280 1235.920 80.540 ;
      LAYER met2 ;
        RECT 589.770 216.650 590.050 220.000 ;
        RECT 589.770 216.510 593.240 216.650 ;
        RECT 589.770 216.000 590.050 216.510 ;
        RECT 593.100 80.570 593.240 216.510 ;
        RECT 593.040 80.250 593.300 80.570 ;
        RECT 1235.660 80.250 1235.920 80.570 ;
        RECT 1235.720 16.730 1235.860 80.250 ;
        RECT 1235.720 16.590 1240.000 16.730 ;
        RECT 1239.860 2.400 1240.000 16.590 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 805.530 1322.500 805.850 1322.560 ;
        RECT 1422.390 1322.500 1422.710 1322.560 ;
        RECT 805.530 1322.360 1422.710 1322.500 ;
        RECT 805.530 1322.300 805.850 1322.360 ;
        RECT 1422.390 1322.300 1422.710 1322.360 ;
        RECT 1257.250 18.600 1257.570 18.660 ;
        RECT 1422.390 18.600 1422.710 18.660 ;
        RECT 1257.250 18.460 1422.710 18.600 ;
        RECT 1257.250 18.400 1257.570 18.460 ;
        RECT 1422.390 18.400 1422.710 18.460 ;
      LAYER via ;
        RECT 805.560 1322.300 805.820 1322.560 ;
        RECT 1422.420 1322.300 1422.680 1322.560 ;
        RECT 1257.280 18.400 1257.540 18.660 ;
        RECT 1422.420 18.400 1422.680 18.660 ;
      LAYER met2 ;
        RECT 804.130 1322.330 804.410 1325.025 ;
        RECT 805.560 1322.330 805.820 1322.590 ;
        RECT 804.130 1322.270 805.820 1322.330 ;
        RECT 1422.420 1322.270 1422.680 1322.590 ;
        RECT 804.130 1322.190 805.760 1322.270 ;
        RECT 804.130 1321.025 804.410 1322.190 ;
        RECT 1422.480 18.690 1422.620 1322.270 ;
        RECT 1257.280 18.370 1257.540 18.690 ;
        RECT 1422.420 18.370 1422.680 18.690 ;
        RECT 1257.340 2.400 1257.480 18.370 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 784.830 1348.340 785.150 1348.400 ;
        RECT 1435.730 1348.340 1436.050 1348.400 ;
        RECT 784.830 1348.200 1436.050 1348.340 ;
        RECT 784.830 1348.140 785.150 1348.200 ;
        RECT 1435.730 1348.140 1436.050 1348.200 ;
        RECT 1275.190 20.640 1275.510 20.700 ;
        RECT 1435.730 20.640 1436.050 20.700 ;
        RECT 1275.190 20.500 1436.050 20.640 ;
        RECT 1275.190 20.440 1275.510 20.500 ;
        RECT 1435.730 20.440 1436.050 20.500 ;
      LAYER via ;
        RECT 784.860 1348.140 785.120 1348.400 ;
        RECT 1435.760 1348.140 1436.020 1348.400 ;
        RECT 1275.220 20.440 1275.480 20.700 ;
        RECT 1435.760 20.440 1436.020 20.700 ;
      LAYER met2 ;
        RECT 784.860 1348.110 785.120 1348.430 ;
        RECT 1435.760 1348.110 1436.020 1348.430 ;
        RECT 784.920 1325.025 785.060 1348.110 ;
        RECT 784.810 1321.025 785.090 1325.025 ;
        RECT 1435.820 20.730 1435.960 1348.110 ;
        RECT 1275.220 20.410 1275.480 20.730 ;
        RECT 1435.760 20.410 1436.020 20.730 ;
        RECT 1275.280 2.400 1275.420 20.410 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1318.045 15.725 1318.215 16.915 ;
      LAYER mcon ;
        RECT 1318.045 16.745 1318.215 16.915 ;
      LAYER met1 ;
        RECT 764.590 1348.000 764.910 1348.060 ;
        RECT 1428.370 1348.000 1428.690 1348.060 ;
        RECT 764.590 1347.860 1428.690 1348.000 ;
        RECT 764.590 1347.800 764.910 1347.860 ;
        RECT 1428.370 1347.800 1428.690 1347.860 ;
        RECT 1317.985 16.900 1318.275 16.945 ;
        RECT 1428.370 16.900 1428.690 16.960 ;
        RECT 1317.985 16.760 1428.690 16.900 ;
        RECT 1317.985 16.715 1318.275 16.760 ;
        RECT 1428.370 16.700 1428.690 16.760 ;
        RECT 1293.130 15.880 1293.450 15.940 ;
        RECT 1317.985 15.880 1318.275 15.925 ;
        RECT 1293.130 15.740 1318.275 15.880 ;
        RECT 1293.130 15.680 1293.450 15.740 ;
        RECT 1317.985 15.695 1318.275 15.740 ;
      LAYER via ;
        RECT 764.620 1347.800 764.880 1348.060 ;
        RECT 1428.400 1347.800 1428.660 1348.060 ;
        RECT 1428.400 16.700 1428.660 16.960 ;
        RECT 1293.160 15.680 1293.420 15.940 ;
      LAYER met2 ;
        RECT 764.620 1347.770 764.880 1348.090 ;
        RECT 1428.400 1347.770 1428.660 1348.090 ;
        RECT 764.680 1325.025 764.820 1347.770 ;
        RECT 764.570 1321.025 764.850 1325.025 ;
        RECT 1428.460 16.990 1428.600 1347.770 ;
        RECT 1428.400 16.670 1428.660 16.990 ;
        RECT 1293.160 15.650 1293.420 15.970 ;
        RECT 1293.220 2.400 1293.360 15.650 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1317.510 197.100 1317.830 197.160 ;
        RECT 1409.970 197.100 1410.290 197.160 ;
        RECT 1317.510 196.960 1410.290 197.100 ;
        RECT 1317.510 196.900 1317.830 196.960 ;
        RECT 1409.970 196.900 1410.290 196.960 ;
        RECT 1311.070 16.900 1311.390 16.960 ;
        RECT 1317.510 16.900 1317.830 16.960 ;
        RECT 1311.070 16.760 1317.830 16.900 ;
        RECT 1311.070 16.700 1311.390 16.760 ;
        RECT 1317.510 16.700 1317.830 16.760 ;
      LAYER via ;
        RECT 1317.540 196.900 1317.800 197.160 ;
        RECT 1410.000 196.900 1410.260 197.160 ;
        RECT 1311.100 16.700 1311.360 16.960 ;
        RECT 1317.540 16.700 1317.800 16.960 ;
      LAYER met2 ;
        RECT 1409.990 929.035 1410.270 929.405 ;
        RECT 1410.060 197.190 1410.200 929.035 ;
        RECT 1317.540 196.870 1317.800 197.190 ;
        RECT 1410.000 196.870 1410.260 197.190 ;
        RECT 1317.600 16.990 1317.740 196.870 ;
        RECT 1311.100 16.670 1311.360 16.990 ;
        RECT 1317.540 16.670 1317.800 16.990 ;
        RECT 1311.160 2.400 1311.300 16.670 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
      LAYER via2 ;
        RECT 1409.990 929.080 1410.270 929.360 ;
      LAYER met3 ;
        RECT 1409.965 929.370 1410.295 929.385 ;
        RECT 1408.060 929.280 1410.295 929.370 ;
        RECT 1404.305 929.070 1410.295 929.280 ;
        RECT 1404.305 928.680 1408.305 929.070 ;
        RECT 1409.965 929.055 1410.295 929.070 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 765.050 142.360 765.370 142.420 ;
        RECT 1324.870 142.360 1325.190 142.420 ;
        RECT 765.050 142.220 1325.190 142.360 ;
        RECT 765.050 142.160 765.370 142.220 ;
        RECT 1324.870 142.160 1325.190 142.220 ;
      LAYER via ;
        RECT 765.080 142.160 765.340 142.420 ;
        RECT 1324.900 142.160 1325.160 142.420 ;
      LAYER met2 ;
        RECT 762.730 216.650 763.010 220.000 ;
        RECT 762.730 216.510 765.280 216.650 ;
        RECT 762.730 216.000 763.010 216.510 ;
        RECT 765.140 142.450 765.280 216.510 ;
        RECT 765.080 142.130 765.340 142.450 ;
        RECT 1324.900 142.130 1325.160 142.450 ;
        RECT 1324.960 17.410 1325.100 142.130 ;
        RECT 1324.960 17.270 1329.240 17.410 ;
        RECT 1329.100 2.400 1329.240 17.270 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 685.085 206.465 685.255 211.055 ;
        RECT 685.085 144.925 685.255 193.035 ;
      LAYER mcon ;
        RECT 685.085 210.885 685.255 211.055 ;
        RECT 685.085 192.865 685.255 193.035 ;
      LAYER met1 ;
        RECT 281.130 1333.720 281.450 1333.780 ;
        RECT 898.910 1333.720 899.230 1333.780 ;
        RECT 281.130 1333.580 899.230 1333.720 ;
        RECT 281.130 1333.520 281.450 1333.580 ;
        RECT 898.910 1333.520 899.230 1333.580 ;
        RECT 281.130 211.040 281.450 211.100 ;
        RECT 685.025 211.040 685.315 211.085 ;
        RECT 281.130 210.900 685.315 211.040 ;
        RECT 281.130 210.840 281.450 210.900 ;
        RECT 685.025 210.855 685.315 210.900 ;
        RECT 685.010 206.620 685.330 206.680 ;
        RECT 684.815 206.480 685.330 206.620 ;
        RECT 685.010 206.420 685.330 206.480 ;
        RECT 685.010 193.020 685.330 193.080 ;
        RECT 684.815 192.880 685.330 193.020 ;
        RECT 685.010 192.820 685.330 192.880 ;
        RECT 685.025 145.080 685.315 145.125 ;
        RECT 685.470 145.080 685.790 145.140 ;
        RECT 685.025 144.940 685.790 145.080 ;
        RECT 685.025 144.895 685.315 144.940 ;
        RECT 685.470 144.880 685.790 144.940 ;
        RECT 683.630 17.240 683.950 17.300 ;
        RECT 686.390 17.240 686.710 17.300 ;
        RECT 683.630 17.100 686.710 17.240 ;
        RECT 683.630 17.040 683.950 17.100 ;
        RECT 686.390 17.040 686.710 17.100 ;
      LAYER via ;
        RECT 281.160 1333.520 281.420 1333.780 ;
        RECT 898.940 1333.520 899.200 1333.780 ;
        RECT 281.160 210.840 281.420 211.100 ;
        RECT 685.040 206.420 685.300 206.680 ;
        RECT 685.040 192.820 685.300 193.080 ;
        RECT 685.500 144.880 685.760 145.140 ;
        RECT 683.660 17.040 683.920 17.300 ;
        RECT 686.420 17.040 686.680 17.300 ;
      LAYER met2 ;
        RECT 281.160 1333.490 281.420 1333.810 ;
        RECT 898.940 1333.490 899.200 1333.810 ;
        RECT 281.220 211.130 281.360 1333.490 ;
        RECT 899.000 1325.025 899.140 1333.490 ;
        RECT 898.890 1321.025 899.170 1325.025 ;
        RECT 281.160 210.810 281.420 211.130 ;
        RECT 685.040 206.390 685.300 206.710 ;
        RECT 685.100 193.110 685.240 206.390 ;
        RECT 685.040 192.790 685.300 193.110 ;
        RECT 685.500 144.850 685.760 145.170 ;
        RECT 685.560 110.570 685.700 144.850 ;
        RECT 684.640 110.430 685.700 110.570 ;
        RECT 684.640 62.290 684.780 110.430 ;
        RECT 683.720 62.150 684.780 62.290 ;
        RECT 683.720 17.330 683.860 62.150 ;
        RECT 683.660 17.010 683.920 17.330 ;
        RECT 686.420 17.010 686.680 17.330 ;
        RECT 686.480 2.400 686.620 17.010 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 836.350 200.500 836.670 200.560 ;
        RECT 840.950 200.500 841.270 200.560 ;
        RECT 836.350 200.360 841.270 200.500 ;
        RECT 836.350 200.300 836.670 200.360 ;
        RECT 840.950 200.300 841.270 200.360 ;
        RECT 840.950 87.620 841.270 87.680 ;
        RECT 1345.570 87.620 1345.890 87.680 ;
        RECT 840.950 87.480 1345.890 87.620 ;
        RECT 840.950 87.420 841.270 87.480 ;
        RECT 1345.570 87.420 1345.890 87.480 ;
      LAYER via ;
        RECT 836.380 200.300 836.640 200.560 ;
        RECT 840.980 200.300 841.240 200.560 ;
        RECT 840.980 87.420 841.240 87.680 ;
        RECT 1345.600 87.420 1345.860 87.680 ;
      LAYER met2 ;
        RECT 836.330 216.000 836.610 220.000 ;
        RECT 836.440 200.590 836.580 216.000 ;
        RECT 836.380 200.270 836.640 200.590 ;
        RECT 840.980 200.270 841.240 200.590 ;
        RECT 841.040 87.710 841.180 200.270 ;
        RECT 840.980 87.390 841.240 87.710 ;
        RECT 1345.600 87.390 1345.860 87.710 ;
        RECT 1345.660 17.410 1345.800 87.390 ;
        RECT 1345.660 17.270 1346.720 17.410 ;
        RECT 1346.580 2.400 1346.720 17.270 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 274.230 1014.460 274.550 1014.520 ;
        RECT 296.770 1014.460 297.090 1014.520 ;
        RECT 274.230 1014.320 297.090 1014.460 ;
        RECT 274.230 1014.260 274.550 1014.320 ;
        RECT 296.770 1014.260 297.090 1014.320 ;
        RECT 274.230 32.880 274.550 32.940 ;
        RECT 1364.430 32.880 1364.750 32.940 ;
        RECT 274.230 32.740 1364.750 32.880 ;
        RECT 274.230 32.680 274.550 32.740 ;
        RECT 1364.430 32.680 1364.750 32.740 ;
      LAYER via ;
        RECT 274.260 1014.260 274.520 1014.520 ;
        RECT 296.800 1014.260 297.060 1014.520 ;
        RECT 274.260 32.680 274.520 32.940 ;
        RECT 1364.460 32.680 1364.720 32.940 ;
      LAYER met2 ;
        RECT 296.790 1016.075 297.070 1016.445 ;
        RECT 296.860 1014.550 297.000 1016.075 ;
        RECT 274.260 1014.230 274.520 1014.550 ;
        RECT 296.800 1014.230 297.060 1014.550 ;
        RECT 274.320 32.970 274.460 1014.230 ;
        RECT 274.260 32.650 274.520 32.970 ;
        RECT 1364.460 32.650 1364.720 32.970 ;
        RECT 1364.520 2.400 1364.660 32.650 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
      LAYER via2 ;
        RECT 296.790 1016.120 297.070 1016.400 ;
      LAYER met3 ;
        RECT 296.765 1016.410 297.095 1016.425 ;
        RECT 296.765 1016.320 310.500 1016.410 ;
        RECT 296.765 1016.110 314.000 1016.320 ;
        RECT 296.765 1016.095 297.095 1016.110 ;
        RECT 310.000 1015.720 314.000 1016.110 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1410.890 638.080 1411.210 638.140 ;
        RECT 1417.790 638.080 1418.110 638.140 ;
        RECT 1410.890 637.940 1418.110 638.080 ;
        RECT 1410.890 637.880 1411.210 637.940 ;
        RECT 1417.790 637.880 1418.110 637.940 ;
        RECT 1407.670 20.300 1407.990 20.360 ;
        RECT 1410.890 20.300 1411.210 20.360 ;
        RECT 1407.670 20.160 1411.210 20.300 ;
        RECT 1407.670 20.100 1407.990 20.160 ;
        RECT 1410.890 20.100 1411.210 20.160 ;
        RECT 1382.370 16.220 1382.690 16.280 ;
        RECT 1407.670 16.220 1407.990 16.280 ;
        RECT 1382.370 16.080 1407.990 16.220 ;
        RECT 1382.370 16.020 1382.690 16.080 ;
        RECT 1407.670 16.020 1407.990 16.080 ;
      LAYER via ;
        RECT 1410.920 637.880 1411.180 638.140 ;
        RECT 1417.820 637.880 1418.080 638.140 ;
        RECT 1407.700 20.100 1407.960 20.360 ;
        RECT 1410.920 20.100 1411.180 20.360 ;
        RECT 1382.400 16.020 1382.660 16.280 ;
        RECT 1407.700 16.020 1407.960 16.280 ;
      LAYER met2 ;
        RECT 1417.810 987.515 1418.090 987.885 ;
        RECT 1417.880 638.170 1418.020 987.515 ;
        RECT 1410.920 637.850 1411.180 638.170 ;
        RECT 1417.820 637.850 1418.080 638.170 ;
        RECT 1410.980 20.390 1411.120 637.850 ;
        RECT 1407.700 20.070 1407.960 20.390 ;
        RECT 1410.920 20.070 1411.180 20.390 ;
        RECT 1407.760 16.310 1407.900 20.070 ;
        RECT 1382.400 15.990 1382.660 16.310 ;
        RECT 1407.700 15.990 1407.960 16.310 ;
        RECT 1382.460 2.400 1382.600 15.990 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
      LAYER via2 ;
        RECT 1417.810 987.560 1418.090 987.840 ;
      LAYER met3 ;
        RECT 1417.785 987.850 1418.115 987.865 ;
        RECT 1408.060 987.760 1418.115 987.850 ;
        RECT 1404.305 987.550 1418.115 987.760 ;
        RECT 1404.305 987.160 1408.305 987.550 ;
        RECT 1417.785 987.535 1418.115 987.550 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 278.370 326.640 278.690 326.700 ;
        RECT 296.770 326.640 297.090 326.700 ;
        RECT 278.370 326.500 297.090 326.640 ;
        RECT 278.370 326.440 278.690 326.500 ;
        RECT 296.770 326.440 297.090 326.500 ;
        RECT 278.370 32.540 278.690 32.600 ;
        RECT 1399.850 32.540 1400.170 32.600 ;
        RECT 278.370 32.400 1400.170 32.540 ;
        RECT 278.370 32.340 278.690 32.400 ;
        RECT 1399.850 32.340 1400.170 32.400 ;
      LAYER via ;
        RECT 278.400 326.440 278.660 326.700 ;
        RECT 296.800 326.440 297.060 326.700 ;
        RECT 278.400 32.340 278.660 32.600 ;
        RECT 1399.880 32.340 1400.140 32.600 ;
      LAYER met2 ;
        RECT 296.790 329.275 297.070 329.645 ;
        RECT 296.860 326.730 297.000 329.275 ;
        RECT 278.400 326.410 278.660 326.730 ;
        RECT 296.800 326.410 297.060 326.730 ;
        RECT 278.460 32.630 278.600 326.410 ;
        RECT 278.400 32.310 278.660 32.630 ;
        RECT 1399.880 32.310 1400.140 32.630 ;
        RECT 1399.940 13.330 1400.080 32.310 ;
        RECT 1399.940 13.190 1400.540 13.330 ;
        RECT 1400.400 2.400 1400.540 13.190 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
      LAYER via2 ;
        RECT 296.790 329.320 297.070 329.600 ;
      LAYER met3 ;
        RECT 296.765 329.610 297.095 329.625 ;
        RECT 296.765 329.520 310.500 329.610 ;
        RECT 296.765 329.310 314.000 329.520 ;
        RECT 296.765 329.295 297.095 329.310 ;
        RECT 310.000 328.920 314.000 329.310 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 910.870 200.500 911.190 200.560 ;
        RECT 916.850 200.500 917.170 200.560 ;
        RECT 910.870 200.360 917.170 200.500 ;
        RECT 910.870 200.300 911.190 200.360 ;
        RECT 916.850 200.300 917.170 200.360 ;
        RECT 916.850 60.080 917.170 60.140 ;
        RECT 1415.030 60.080 1415.350 60.140 ;
        RECT 916.850 59.940 1415.350 60.080 ;
        RECT 916.850 59.880 917.170 59.940 ;
        RECT 1415.030 59.880 1415.350 59.940 ;
      LAYER via ;
        RECT 910.900 200.300 911.160 200.560 ;
        RECT 916.880 200.300 917.140 200.560 ;
        RECT 916.880 59.880 917.140 60.140 ;
        RECT 1415.060 59.880 1415.320 60.140 ;
      LAYER met2 ;
        RECT 910.850 216.000 911.130 220.000 ;
        RECT 910.960 200.590 911.100 216.000 ;
        RECT 910.900 200.270 911.160 200.590 ;
        RECT 916.880 200.270 917.140 200.590 ;
        RECT 916.940 60.170 917.080 200.270 ;
        RECT 916.880 59.850 917.140 60.170 ;
        RECT 1415.060 59.850 1415.320 60.170 ;
        RECT 1415.120 16.900 1415.260 59.850 ;
        RECT 1415.120 16.760 1418.480 16.900 ;
        RECT 1418.340 2.400 1418.480 16.760 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1395.710 200.500 1396.030 200.560 ;
        RECT 1400.310 200.500 1400.630 200.560 ;
        RECT 1395.710 200.360 1400.630 200.500 ;
        RECT 1395.710 200.300 1396.030 200.360 ;
        RECT 1400.310 200.300 1400.630 200.360 ;
        RECT 1400.310 156.640 1400.630 156.700 ;
        RECT 1436.190 156.640 1436.510 156.700 ;
        RECT 1400.310 156.500 1436.510 156.640 ;
        RECT 1400.310 156.440 1400.630 156.500 ;
        RECT 1436.190 156.440 1436.510 156.500 ;
      LAYER via ;
        RECT 1395.740 200.300 1396.000 200.560 ;
        RECT 1400.340 200.300 1400.600 200.560 ;
        RECT 1400.340 156.440 1400.600 156.700 ;
        RECT 1436.220 156.440 1436.480 156.700 ;
      LAYER met2 ;
        RECT 1395.690 216.000 1395.970 220.000 ;
        RECT 1395.800 200.590 1395.940 216.000 ;
        RECT 1395.740 200.270 1396.000 200.590 ;
        RECT 1400.340 200.270 1400.600 200.590 ;
        RECT 1400.400 156.730 1400.540 200.270 ;
        RECT 1400.340 156.410 1400.600 156.730 ;
        RECT 1436.220 156.410 1436.480 156.730 ;
        RECT 1436.280 17.410 1436.420 156.410 ;
        RECT 1435.820 17.270 1436.420 17.410 ;
        RECT 1435.820 2.400 1435.960 17.270 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 317.800 1419.490 317.860 ;
        RECT 1449.530 317.800 1449.850 317.860 ;
        RECT 1419.170 317.660 1449.850 317.800 ;
        RECT 1419.170 317.600 1419.490 317.660 ;
        RECT 1449.530 317.600 1449.850 317.660 ;
      LAYER via ;
        RECT 1419.200 317.600 1419.460 317.860 ;
        RECT 1449.560 317.600 1449.820 317.860 ;
      LAYER met2 ;
        RECT 1419.190 322.475 1419.470 322.845 ;
        RECT 1419.260 317.890 1419.400 322.475 ;
        RECT 1419.200 317.570 1419.460 317.890 ;
        RECT 1449.560 317.570 1449.820 317.890 ;
        RECT 1449.620 16.730 1449.760 317.570 ;
        RECT 1449.620 16.590 1453.900 16.730 ;
        RECT 1453.760 2.400 1453.900 16.590 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
      LAYER via2 ;
        RECT 1419.190 322.520 1419.470 322.800 ;
      LAYER met3 ;
        RECT 1419.165 322.810 1419.495 322.825 ;
        RECT 1408.060 322.720 1419.495 322.810 ;
        RECT 1404.305 322.510 1419.495 322.720 ;
        RECT 1404.305 322.120 1408.305 322.510 ;
        RECT 1419.165 322.495 1419.495 322.510 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 265.950 904.300 266.270 904.360 ;
        RECT 296.770 904.300 297.090 904.360 ;
        RECT 265.950 904.160 297.090 904.300 ;
        RECT 265.950 904.100 266.270 904.160 ;
        RECT 296.770 904.100 297.090 904.160 ;
        RECT 265.950 45.800 266.270 45.860 ;
        RECT 1471.610 45.800 1471.930 45.860 ;
        RECT 265.950 45.660 1471.930 45.800 ;
        RECT 265.950 45.600 266.270 45.660 ;
        RECT 1471.610 45.600 1471.930 45.660 ;
      LAYER via ;
        RECT 265.980 904.100 266.240 904.360 ;
        RECT 296.800 904.100 297.060 904.360 ;
        RECT 265.980 45.600 266.240 45.860 ;
        RECT 1471.640 45.600 1471.900 45.860 ;
      LAYER met2 ;
        RECT 296.790 907.275 297.070 907.645 ;
        RECT 296.860 904.390 297.000 907.275 ;
        RECT 265.980 904.070 266.240 904.390 ;
        RECT 296.800 904.070 297.060 904.390 ;
        RECT 266.040 45.890 266.180 904.070 ;
        RECT 265.980 45.570 266.240 45.890 ;
        RECT 1471.640 45.570 1471.900 45.890 ;
        RECT 1471.700 2.400 1471.840 45.570 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
      LAYER via2 ;
        RECT 296.790 907.320 297.070 907.600 ;
      LAYER met3 ;
        RECT 296.765 907.610 297.095 907.625 ;
        RECT 296.765 907.520 310.500 907.610 ;
        RECT 296.765 907.310 314.000 907.520 ;
        RECT 296.765 907.295 297.095 907.310 ;
        RECT 310.000 906.920 314.000 907.310 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 682.250 1321.820 682.570 1321.880 ;
        RECT 682.250 1321.680 722.500 1321.820 ;
        RECT 682.250 1321.620 682.570 1321.680 ;
        RECT 722.360 1320.800 722.500 1321.680 ;
        RECT 1483.570 1320.800 1483.890 1320.860 ;
        RECT 722.360 1320.660 1483.890 1320.800 ;
        RECT 1483.570 1320.600 1483.890 1320.660 ;
        RECT 1483.570 16.900 1483.890 16.960 ;
        RECT 1489.550 16.900 1489.870 16.960 ;
        RECT 1483.570 16.760 1489.870 16.900 ;
        RECT 1483.570 16.700 1483.890 16.760 ;
        RECT 1489.550 16.700 1489.870 16.760 ;
      LAYER via ;
        RECT 682.280 1321.620 682.540 1321.880 ;
        RECT 1483.600 1320.600 1483.860 1320.860 ;
        RECT 1483.600 16.700 1483.860 16.960 ;
        RECT 1489.580 16.700 1489.840 16.960 ;
      LAYER met2 ;
        RECT 680.850 1321.650 681.130 1325.025 ;
        RECT 682.280 1321.650 682.540 1321.910 ;
        RECT 680.850 1321.590 682.540 1321.650 ;
        RECT 680.850 1321.510 682.480 1321.590 ;
        RECT 680.850 1321.025 681.130 1321.510 ;
        RECT 1483.600 1320.570 1483.860 1320.890 ;
        RECT 1483.660 16.990 1483.800 1320.570 ;
        RECT 1483.600 16.670 1483.860 16.990 ;
        RECT 1489.580 16.670 1489.840 16.990 ;
        RECT 1489.640 2.400 1489.780 16.670 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1211.250 1321.820 1211.570 1321.880 ;
        RECT 1504.270 1321.820 1504.590 1321.880 ;
        RECT 1211.250 1321.680 1504.590 1321.820 ;
        RECT 1211.250 1321.620 1211.570 1321.680 ;
        RECT 1504.270 1321.620 1504.590 1321.680 ;
      LAYER via ;
        RECT 1211.280 1321.620 1211.540 1321.880 ;
        RECT 1504.300 1321.620 1504.560 1321.880 ;
      LAYER met2 ;
        RECT 1209.850 1321.650 1210.130 1325.025 ;
        RECT 1211.280 1321.650 1211.540 1321.910 ;
        RECT 1209.850 1321.590 1211.540 1321.650 ;
        RECT 1504.300 1321.590 1504.560 1321.910 ;
        RECT 1209.850 1321.510 1211.480 1321.590 ;
        RECT 1209.850 1321.025 1210.130 1321.510 ;
        RECT 1504.360 17.410 1504.500 1321.590 ;
        RECT 1504.360 17.270 1507.260 17.410 ;
        RECT 1507.120 2.400 1507.260 17.270 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 704.330 17.240 704.650 17.300 ;
        RECT 710.310 17.240 710.630 17.300 ;
        RECT 704.330 17.100 710.630 17.240 ;
        RECT 704.330 17.040 704.650 17.100 ;
        RECT 710.310 17.040 710.630 17.100 ;
      LAYER via ;
        RECT 704.360 17.040 704.620 17.300 ;
        RECT 710.340 17.040 710.600 17.300 ;
      LAYER met2 ;
        RECT 1001.970 1339.755 1002.250 1340.125 ;
        RECT 1002.040 1325.025 1002.180 1339.755 ;
        RECT 1001.930 1321.025 1002.210 1325.025 ;
        RECT 710.330 217.075 710.610 217.445 ;
        RECT 710.400 17.330 710.540 217.075 ;
        RECT 704.360 17.010 704.620 17.330 ;
        RECT 710.340 17.010 710.600 17.330 ;
        RECT 704.420 2.400 704.560 17.010 ;
        RECT 704.210 -4.800 704.770 2.400 ;
      LAYER via2 ;
        RECT 1001.970 1339.800 1002.250 1340.080 ;
        RECT 710.330 217.120 710.610 217.400 ;
      LAYER met3 ;
        RECT 1001.945 1340.090 1002.275 1340.105 ;
        RECT 1408.790 1340.090 1409.170 1340.100 ;
        RECT 1001.945 1339.790 1409.170 1340.090 ;
        RECT 1001.945 1339.775 1002.275 1339.790 ;
        RECT 1408.790 1339.780 1409.170 1339.790 ;
        RECT 710.305 217.410 710.635 217.425 ;
        RECT 1408.790 217.410 1409.170 217.420 ;
        RECT 710.305 217.110 1409.170 217.410 ;
        RECT 710.305 217.095 710.635 217.110 ;
        RECT 1408.790 217.100 1409.170 217.110 ;
      LAYER via3 ;
        RECT 1408.820 1339.780 1409.140 1340.100 ;
        RECT 1408.820 217.100 1409.140 217.420 ;
      LAYER met4 ;
        RECT 1408.815 1339.775 1409.145 1340.105 ;
        RECT 1408.830 217.425 1409.130 1339.775 ;
        RECT 1408.815 217.095 1409.145 217.425 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 423.270 1335.420 423.590 1335.480 ;
        RECT 1524.970 1335.420 1525.290 1335.480 ;
        RECT 423.270 1335.280 1525.290 1335.420 ;
        RECT 423.270 1335.220 423.590 1335.280 ;
        RECT 1524.970 1335.220 1525.290 1335.280 ;
      LAYER via ;
        RECT 423.300 1335.220 423.560 1335.480 ;
        RECT 1525.000 1335.220 1525.260 1335.480 ;
      LAYER met2 ;
        RECT 423.300 1335.190 423.560 1335.510 ;
        RECT 1525.000 1335.190 1525.260 1335.510 ;
        RECT 423.360 1325.025 423.500 1335.190 ;
        RECT 423.250 1321.025 423.530 1325.025 ;
        RECT 1525.060 2.400 1525.200 1335.190 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.390 200.500 594.710 200.560 ;
        RECT 599.450 200.500 599.770 200.560 ;
        RECT 594.390 200.360 599.770 200.500 ;
        RECT 594.390 200.300 594.710 200.360 ;
        RECT 599.450 200.300 599.770 200.360 ;
        RECT 599.450 156.300 599.770 156.360 ;
        RECT 1538.770 156.300 1539.090 156.360 ;
        RECT 599.450 156.160 1539.090 156.300 ;
        RECT 599.450 156.100 599.770 156.160 ;
        RECT 1538.770 156.100 1539.090 156.160 ;
      LAYER via ;
        RECT 594.420 200.300 594.680 200.560 ;
        RECT 599.480 200.300 599.740 200.560 ;
        RECT 599.480 156.100 599.740 156.360 ;
        RECT 1538.800 156.100 1539.060 156.360 ;
      LAYER met2 ;
        RECT 594.370 216.000 594.650 220.000 ;
        RECT 594.480 200.590 594.620 216.000 ;
        RECT 594.420 200.270 594.680 200.590 ;
        RECT 599.480 200.270 599.740 200.590 ;
        RECT 599.540 156.390 599.680 200.270 ;
        RECT 599.480 156.070 599.740 156.390 ;
        RECT 1538.800 156.070 1539.060 156.390 ;
        RECT 1538.860 17.410 1539.000 156.070 ;
        RECT 1538.860 17.270 1543.140 17.410 ;
        RECT 1543.000 2.400 1543.140 17.270 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1228.320 1421.330 1228.380 ;
        RECT 1559.470 1228.320 1559.790 1228.380 ;
        RECT 1421.010 1228.180 1559.790 1228.320 ;
        RECT 1421.010 1228.120 1421.330 1228.180 ;
        RECT 1559.470 1228.120 1559.790 1228.180 ;
      LAYER via ;
        RECT 1421.040 1228.120 1421.300 1228.380 ;
        RECT 1559.500 1228.120 1559.760 1228.380 ;
      LAYER met2 ;
        RECT 1421.030 1228.235 1421.310 1228.605 ;
        RECT 1421.040 1228.090 1421.300 1228.235 ;
        RECT 1559.500 1228.090 1559.760 1228.410 ;
        RECT 1559.560 17.410 1559.700 1228.090 ;
        RECT 1559.560 17.270 1561.080 17.410 ;
        RECT 1560.940 2.400 1561.080 17.270 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1228.280 1421.310 1228.560 ;
      LAYER met3 ;
        RECT 1421.005 1228.570 1421.335 1228.585 ;
        RECT 1408.060 1228.480 1421.335 1228.570 ;
        RECT 1404.305 1228.270 1421.335 1228.480 ;
        RECT 1404.305 1227.880 1408.305 1228.270 ;
        RECT 1421.005 1228.255 1421.335 1228.270 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 273.310 600.680 273.630 600.740 ;
        RECT 296.770 600.680 297.090 600.740 ;
        RECT 273.310 600.540 297.090 600.680 ;
        RECT 273.310 600.480 273.630 600.540 ;
        RECT 296.770 600.480 297.090 600.540 ;
        RECT 273.310 45.460 273.630 45.520 ;
        RECT 1578.790 45.460 1579.110 45.520 ;
        RECT 273.310 45.320 1579.110 45.460 ;
        RECT 273.310 45.260 273.630 45.320 ;
        RECT 1578.790 45.260 1579.110 45.320 ;
      LAYER via ;
        RECT 273.340 600.480 273.600 600.740 ;
        RECT 296.800 600.480 297.060 600.740 ;
        RECT 273.340 45.260 273.600 45.520 ;
        RECT 1578.820 45.260 1579.080 45.520 ;
      LAYER met2 ;
        RECT 296.790 606.715 297.070 607.085 ;
        RECT 296.860 600.770 297.000 606.715 ;
        RECT 273.340 600.450 273.600 600.770 ;
        RECT 296.800 600.450 297.060 600.770 ;
        RECT 273.400 45.550 273.540 600.450 ;
        RECT 273.340 45.230 273.600 45.550 ;
        RECT 1578.820 45.230 1579.080 45.550 ;
        RECT 1578.880 2.400 1579.020 45.230 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
      LAYER via2 ;
        RECT 296.790 606.760 297.070 607.040 ;
      LAYER met3 ;
        RECT 296.765 607.050 297.095 607.065 ;
        RECT 296.765 606.960 310.500 607.050 ;
        RECT 296.765 606.750 314.000 606.960 ;
        RECT 296.765 606.735 297.095 606.750 ;
        RECT 310.000 606.360 314.000 606.750 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 744.350 121.620 744.670 121.680 ;
        RECT 1593.970 121.620 1594.290 121.680 ;
        RECT 744.350 121.480 1594.290 121.620 ;
        RECT 744.350 121.420 744.670 121.480 ;
        RECT 1593.970 121.420 1594.290 121.480 ;
        RECT 1593.970 2.960 1594.290 3.020 ;
        RECT 1596.270 2.960 1596.590 3.020 ;
        RECT 1593.970 2.820 1596.590 2.960 ;
        RECT 1593.970 2.760 1594.290 2.820 ;
        RECT 1596.270 2.760 1596.590 2.820 ;
      LAYER via ;
        RECT 744.380 121.420 744.640 121.680 ;
        RECT 1594.000 121.420 1594.260 121.680 ;
        RECT 1594.000 2.760 1594.260 3.020 ;
        RECT 1596.300 2.760 1596.560 3.020 ;
      LAYER met2 ;
        RECT 742.490 216.650 742.770 220.000 ;
        RECT 742.490 216.510 744.580 216.650 ;
        RECT 742.490 216.000 742.770 216.510 ;
        RECT 744.440 121.710 744.580 216.510 ;
        RECT 744.380 121.390 744.640 121.710 ;
        RECT 1594.000 121.390 1594.260 121.710 ;
        RECT 1594.060 3.050 1594.200 121.390 ;
        RECT 1594.000 2.730 1594.260 3.050 ;
        RECT 1596.300 2.730 1596.560 3.050 ;
        RECT 1596.360 2.400 1596.500 2.730 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1048.870 200.500 1049.190 200.560 ;
        RECT 1054.850 200.500 1055.170 200.560 ;
        RECT 1048.870 200.360 1055.170 200.500 ;
        RECT 1048.870 200.300 1049.190 200.360 ;
        RECT 1054.850 200.300 1055.170 200.360 ;
        RECT 1054.850 73.340 1055.170 73.400 ;
        RECT 1607.770 73.340 1608.090 73.400 ;
        RECT 1054.850 73.200 1608.090 73.340 ;
        RECT 1054.850 73.140 1055.170 73.200 ;
        RECT 1607.770 73.140 1608.090 73.200 ;
        RECT 1607.770 16.900 1608.090 16.960 ;
        RECT 1614.210 16.900 1614.530 16.960 ;
        RECT 1607.770 16.760 1614.530 16.900 ;
        RECT 1607.770 16.700 1608.090 16.760 ;
        RECT 1614.210 16.700 1614.530 16.760 ;
      LAYER via ;
        RECT 1048.900 200.300 1049.160 200.560 ;
        RECT 1054.880 200.300 1055.140 200.560 ;
        RECT 1054.880 73.140 1055.140 73.400 ;
        RECT 1607.800 73.140 1608.060 73.400 ;
        RECT 1607.800 16.700 1608.060 16.960 ;
        RECT 1614.240 16.700 1614.500 16.960 ;
      LAYER met2 ;
        RECT 1048.850 216.000 1049.130 220.000 ;
        RECT 1048.960 200.590 1049.100 216.000 ;
        RECT 1048.900 200.270 1049.160 200.590 ;
        RECT 1054.880 200.270 1055.140 200.590 ;
        RECT 1054.940 73.430 1055.080 200.270 ;
        RECT 1054.880 73.110 1055.140 73.430 ;
        RECT 1607.800 73.110 1608.060 73.430 ;
        RECT 1607.860 16.990 1608.000 73.110 ;
        RECT 1607.800 16.670 1608.060 16.990 ;
        RECT 1614.240 16.670 1614.500 16.990 ;
        RECT 1614.300 2.400 1614.440 16.670 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 266.410 966.180 266.730 966.240 ;
        RECT 296.770 966.180 297.090 966.240 ;
        RECT 266.410 966.040 297.090 966.180 ;
        RECT 266.410 965.980 266.730 966.040 ;
        RECT 296.770 965.980 297.090 966.040 ;
        RECT 266.410 45.120 266.730 45.180 ;
        RECT 1632.150 45.120 1632.470 45.180 ;
        RECT 266.410 44.980 1632.470 45.120 ;
        RECT 266.410 44.920 266.730 44.980 ;
        RECT 1632.150 44.920 1632.470 44.980 ;
      LAYER via ;
        RECT 266.440 965.980 266.700 966.240 ;
        RECT 296.800 965.980 297.060 966.240 ;
        RECT 266.440 44.920 266.700 45.180 ;
        RECT 1632.180 44.920 1632.440 45.180 ;
      LAYER met2 ;
        RECT 296.790 972.555 297.070 972.925 ;
        RECT 296.860 966.270 297.000 972.555 ;
        RECT 266.440 965.950 266.700 966.270 ;
        RECT 296.800 965.950 297.060 966.270 ;
        RECT 266.500 45.210 266.640 965.950 ;
        RECT 266.440 44.890 266.700 45.210 ;
        RECT 1632.180 44.890 1632.440 45.210 ;
        RECT 1632.240 2.400 1632.380 44.890 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
      LAYER via2 ;
        RECT 296.790 972.600 297.070 972.880 ;
      LAYER met3 ;
        RECT 296.765 972.890 297.095 972.905 ;
        RECT 296.765 972.800 310.500 972.890 ;
        RECT 296.765 972.590 314.000 972.800 ;
        RECT 296.765 972.575 297.095 972.590 ;
        RECT 310.000 972.200 314.000 972.590 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.610 1321.650 1373.890 1325.025 ;
        RECT 1375.030 1321.650 1375.310 1321.765 ;
        RECT 1373.610 1321.510 1375.310 1321.650 ;
        RECT 1373.610 1321.025 1373.890 1321.510 ;
        RECT 1375.030 1321.395 1375.310 1321.510 ;
        RECT 1650.110 15.795 1650.390 16.165 ;
        RECT 1650.180 2.400 1650.320 15.795 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
      LAYER via2 ;
        RECT 1375.030 1321.440 1375.310 1321.720 ;
        RECT 1650.110 15.840 1650.390 16.120 ;
      LAYER met3 ;
        RECT 1375.005 1321.730 1375.335 1321.745 ;
        RECT 1396.830 1321.730 1397.210 1321.740 ;
        RECT 1375.005 1321.430 1397.210 1321.730 ;
        RECT 1375.005 1321.415 1375.335 1321.430 ;
        RECT 1396.830 1321.420 1397.210 1321.430 ;
        RECT 1396.830 16.130 1397.210 16.140 ;
        RECT 1650.085 16.130 1650.415 16.145 ;
        RECT 1396.830 15.830 1650.415 16.130 ;
        RECT 1396.830 15.820 1397.210 15.830 ;
        RECT 1650.085 15.815 1650.415 15.830 ;
      LAYER via3 ;
        RECT 1396.860 1321.420 1397.180 1321.740 ;
        RECT 1396.860 15.820 1397.180 16.140 ;
      LAYER met4 ;
        RECT 1396.855 1321.415 1397.185 1321.745 ;
        RECT 1396.870 16.145 1397.170 1321.415 ;
        RECT 1396.855 15.815 1397.185 16.145 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1420.550 1256.200 1420.870 1256.260 ;
        RECT 1662.970 1256.200 1663.290 1256.260 ;
        RECT 1420.550 1256.060 1663.290 1256.200 ;
        RECT 1420.550 1256.000 1420.870 1256.060 ;
        RECT 1662.970 1256.000 1663.290 1256.060 ;
      LAYER via ;
        RECT 1420.580 1256.000 1420.840 1256.260 ;
        RECT 1663.000 1256.000 1663.260 1256.260 ;
      LAYER met2 ;
        RECT 1420.570 1258.155 1420.850 1258.525 ;
        RECT 1420.640 1256.290 1420.780 1258.155 ;
        RECT 1420.580 1255.970 1420.840 1256.290 ;
        RECT 1663.000 1255.970 1663.260 1256.290 ;
        RECT 1663.060 17.410 1663.200 1255.970 ;
        RECT 1663.060 17.270 1668.260 17.410 ;
        RECT 1668.120 2.400 1668.260 17.270 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
      LAYER via2 ;
        RECT 1420.570 1258.200 1420.850 1258.480 ;
      LAYER met3 ;
        RECT 1420.545 1258.490 1420.875 1258.505 ;
        RECT 1408.060 1258.400 1420.875 1258.490 ;
        RECT 1404.305 1258.190 1420.875 1258.400 ;
        RECT 1404.305 1257.800 1408.305 1258.190 ;
        RECT 1420.545 1258.175 1420.875 1258.190 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 654.650 114.480 654.970 114.540 ;
        RECT 1683.670 114.480 1683.990 114.540 ;
        RECT 654.650 114.340 1683.990 114.480 ;
        RECT 654.650 114.280 654.970 114.340 ;
        RECT 1683.670 114.280 1683.990 114.340 ;
      LAYER via ;
        RECT 654.680 114.280 654.940 114.540 ;
        RECT 1683.700 114.280 1683.960 114.540 ;
      LAYER met2 ;
        RECT 653.250 216.650 653.530 220.000 ;
        RECT 653.250 216.510 654.880 216.650 ;
        RECT 653.250 216.000 653.530 216.510 ;
        RECT 654.740 114.570 654.880 216.510 ;
        RECT 654.680 114.250 654.940 114.570 ;
        RECT 1683.700 114.250 1683.960 114.570 ;
        RECT 1683.760 17.410 1683.900 114.250 ;
        RECT 1683.760 17.270 1685.740 17.410 ;
        RECT 1685.600 2.400 1685.740 17.270 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 722.270 33.560 722.590 33.620 ;
        RECT 1118.330 33.560 1118.650 33.620 ;
        RECT 722.270 33.420 1118.650 33.560 ;
        RECT 722.270 33.360 722.590 33.420 ;
        RECT 1118.330 33.360 1118.650 33.420 ;
      LAYER via ;
        RECT 722.300 33.360 722.560 33.620 ;
        RECT 1118.360 33.360 1118.620 33.620 ;
      LAYER met2 ;
        RECT 1118.770 216.650 1119.050 220.000 ;
        RECT 1118.420 216.510 1119.050 216.650 ;
        RECT 1118.420 33.650 1118.560 216.510 ;
        RECT 1118.770 216.000 1119.050 216.510 ;
        RECT 722.300 33.330 722.560 33.650 ;
        RECT 1118.360 33.330 1118.620 33.650 ;
        RECT 722.360 2.400 722.500 33.330 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.410 1321.650 1111.690 1325.025 ;
        RECT 1112.830 1321.650 1113.110 1321.765 ;
        RECT 1111.410 1321.510 1113.110 1321.650 ;
        RECT 1111.410 1321.025 1111.690 1321.510 ;
        RECT 1112.830 1321.395 1113.110 1321.510 ;
        RECT 1703.470 19.875 1703.750 20.245 ;
        RECT 1703.540 2.400 1703.680 19.875 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
      LAYER via2 ;
        RECT 1112.830 1321.440 1113.110 1321.720 ;
        RECT 1703.470 19.920 1703.750 20.200 ;
      LAYER met3 ;
        RECT 1112.805 1321.730 1113.135 1321.745 ;
        RECT 1124.510 1321.730 1124.890 1321.740 ;
        RECT 1112.805 1321.430 1124.890 1321.730 ;
        RECT 1112.805 1321.415 1113.135 1321.430 ;
        RECT 1124.510 1321.420 1124.890 1321.430 ;
        RECT 1124.510 1320.370 1124.890 1320.380 ;
        RECT 1405.110 1320.370 1405.490 1320.380 ;
        RECT 1124.510 1320.070 1405.490 1320.370 ;
        RECT 1124.510 1320.060 1124.890 1320.070 ;
        RECT 1405.110 1320.060 1405.490 1320.070 ;
        RECT 1405.110 20.210 1405.490 20.220 ;
        RECT 1703.445 20.210 1703.775 20.225 ;
        RECT 1405.110 19.910 1703.775 20.210 ;
        RECT 1405.110 19.900 1405.490 19.910 ;
        RECT 1703.445 19.895 1703.775 19.910 ;
      LAYER via3 ;
        RECT 1124.540 1321.420 1124.860 1321.740 ;
        RECT 1124.540 1320.060 1124.860 1320.380 ;
        RECT 1405.140 1320.060 1405.460 1320.380 ;
        RECT 1405.140 19.900 1405.460 20.220 ;
      LAYER met4 ;
        RECT 1124.535 1321.415 1124.865 1321.745 ;
        RECT 1124.550 1320.385 1124.850 1321.415 ;
        RECT 1124.535 1320.055 1124.865 1320.385 ;
        RECT 1405.135 1320.055 1405.465 1320.385 ;
        RECT 1405.150 20.225 1405.450 1320.055 ;
        RECT 1405.135 19.895 1405.465 20.225 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 945.830 200.500 946.150 200.560 ;
        RECT 951.810 200.500 952.130 200.560 ;
        RECT 945.830 200.360 952.130 200.500 ;
        RECT 945.830 200.300 946.150 200.360 ;
        RECT 951.810 200.300 952.130 200.360 ;
        RECT 951.810 65.860 952.130 65.920 ;
        RECT 1718.170 65.860 1718.490 65.920 ;
        RECT 951.810 65.720 1718.490 65.860 ;
        RECT 951.810 65.660 952.130 65.720 ;
        RECT 1718.170 65.660 1718.490 65.720 ;
      LAYER via ;
        RECT 945.860 200.300 946.120 200.560 ;
        RECT 951.840 200.300 952.100 200.560 ;
        RECT 951.840 65.660 952.100 65.920 ;
        RECT 1718.200 65.660 1718.460 65.920 ;
      LAYER met2 ;
        RECT 945.810 216.000 946.090 220.000 ;
        RECT 945.920 200.590 946.060 216.000 ;
        RECT 945.860 200.270 946.120 200.590 ;
        RECT 951.840 200.270 952.100 200.590 ;
        RECT 951.900 65.950 952.040 200.270 ;
        RECT 951.840 65.630 952.100 65.950 ;
        RECT 1718.200 65.630 1718.460 65.950 ;
        RECT 1718.260 17.410 1718.400 65.630 ;
        RECT 1718.260 17.270 1721.620 17.410 ;
        RECT 1721.480 2.400 1721.620 17.270 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1418.250 586.740 1418.570 586.800 ;
        RECT 1739.330 586.740 1739.650 586.800 ;
        RECT 1418.250 586.600 1739.650 586.740 ;
        RECT 1418.250 586.540 1418.570 586.600 ;
        RECT 1739.330 586.540 1739.650 586.600 ;
      LAYER via ;
        RECT 1418.280 586.540 1418.540 586.800 ;
        RECT 1739.360 586.540 1739.620 586.800 ;
      LAYER met2 ;
        RECT 1418.270 593.115 1418.550 593.485 ;
        RECT 1418.340 586.830 1418.480 593.115 ;
        RECT 1418.280 586.510 1418.540 586.830 ;
        RECT 1739.360 586.510 1739.620 586.830 ;
        RECT 1739.420 2.400 1739.560 586.510 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
      LAYER via2 ;
        RECT 1418.270 593.160 1418.550 593.440 ;
      LAYER met3 ;
        RECT 1418.245 593.450 1418.575 593.465 ;
        RECT 1408.060 593.360 1418.575 593.450 ;
        RECT 1404.305 593.150 1418.575 593.360 ;
        RECT 1404.305 592.760 1408.305 593.150 ;
        RECT 1418.245 593.135 1418.575 593.150 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 302.750 142.020 303.070 142.080 ;
        RECT 1752.670 142.020 1752.990 142.080 ;
        RECT 302.750 141.880 1752.990 142.020 ;
        RECT 302.750 141.820 303.070 141.880 ;
        RECT 1752.670 141.820 1752.990 141.880 ;
      LAYER via ;
        RECT 302.780 141.820 303.040 142.080 ;
        RECT 1752.700 141.820 1752.960 142.080 ;
      LAYER met2 ;
        RECT 306.910 489.755 307.190 490.125 ;
        RECT 306.980 488.765 307.120 489.755 ;
        RECT 302.770 488.395 303.050 488.765 ;
        RECT 306.910 488.395 307.190 488.765 ;
        RECT 302.840 142.110 302.980 488.395 ;
        RECT 302.780 141.790 303.040 142.110 ;
        RECT 1752.700 141.790 1752.960 142.110 ;
        RECT 1752.760 17.410 1752.900 141.790 ;
        RECT 1752.760 17.270 1757.040 17.410 ;
        RECT 1756.900 2.400 1757.040 17.270 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
      LAYER via2 ;
        RECT 306.910 489.800 307.190 490.080 ;
        RECT 302.770 488.440 303.050 488.720 ;
        RECT 306.910 488.440 307.190 488.720 ;
      LAYER met3 ;
        RECT 306.885 490.090 307.215 490.105 ;
        RECT 302.990 489.790 307.215 490.090 ;
        RECT 302.990 488.745 303.290 489.790 ;
        RECT 306.885 489.775 307.215 489.790 ;
        RECT 310.000 489.400 314.000 490.000 ;
        RECT 302.745 488.430 303.290 488.745 ;
        RECT 306.885 488.730 307.215 488.745 ;
        RECT 311.270 488.730 311.570 489.400 ;
        RECT 306.885 488.430 311.570 488.730 ;
        RECT 302.745 488.415 303.075 488.430 ;
        RECT 306.885 488.415 307.215 488.430 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 676.500 1421.330 676.560 ;
        RECT 1773.370 676.500 1773.690 676.560 ;
        RECT 1421.010 676.360 1773.690 676.500 ;
        RECT 1421.010 676.300 1421.330 676.360 ;
        RECT 1773.370 676.300 1773.690 676.360 ;
      LAYER via ;
        RECT 1421.040 676.300 1421.300 676.560 ;
        RECT 1773.400 676.300 1773.660 676.560 ;
      LAYER met2 ;
        RECT 1421.030 680.155 1421.310 680.525 ;
        RECT 1421.100 676.590 1421.240 680.155 ;
        RECT 1421.040 676.270 1421.300 676.590 ;
        RECT 1773.400 676.270 1773.660 676.590 ;
        RECT 1773.460 17.410 1773.600 676.270 ;
        RECT 1773.460 17.270 1774.980 17.410 ;
        RECT 1774.840 2.400 1774.980 17.270 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
      LAYER via2 ;
        RECT 1421.030 680.200 1421.310 680.480 ;
      LAYER met3 ;
        RECT 1421.005 680.490 1421.335 680.505 ;
        RECT 1408.060 680.400 1421.335 680.490 ;
        RECT 1404.305 680.190 1421.335 680.400 ;
        RECT 1404.305 679.800 1408.305 680.190 ;
        RECT 1421.005 680.175 1421.335 680.190 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1122.085 1314.525 1122.255 1321.495 ;
      LAYER mcon ;
        RECT 1122.085 1321.325 1122.255 1321.495 ;
      LAYER met1 ;
        RECT 1122.010 1321.480 1122.330 1321.540 ;
        RECT 1121.815 1321.340 1122.330 1321.480 ;
        RECT 1122.010 1321.280 1122.330 1321.340 ;
        RECT 1122.025 1314.680 1122.315 1314.725 ;
        RECT 1787.170 1314.680 1787.490 1314.740 ;
        RECT 1122.025 1314.540 1787.490 1314.680 ;
        RECT 1122.025 1314.495 1122.315 1314.540 ;
        RECT 1787.170 1314.480 1787.490 1314.540 ;
      LAYER via ;
        RECT 1122.040 1321.280 1122.300 1321.540 ;
        RECT 1787.200 1314.480 1787.460 1314.740 ;
      LAYER met2 ;
        RECT 1120.610 1321.650 1120.890 1325.025 ;
        RECT 1120.610 1321.570 1122.240 1321.650 ;
        RECT 1120.610 1321.510 1122.300 1321.570 ;
        RECT 1120.610 1321.025 1120.890 1321.510 ;
        RECT 1122.040 1321.250 1122.300 1321.510 ;
        RECT 1787.200 1314.450 1787.460 1314.770 ;
        RECT 1787.260 17.410 1787.400 1314.450 ;
        RECT 1787.260 17.270 1792.920 17.410 ;
        RECT 1792.780 2.400 1792.920 17.270 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 661.550 1321.280 661.870 1321.540 ;
        RECT 661.640 1319.780 661.780 1321.280 ;
        RECT 1807.870 1319.780 1808.190 1319.840 ;
        RECT 661.640 1319.640 1808.190 1319.780 ;
        RECT 1807.870 1319.580 1808.190 1319.640 ;
      LAYER via ;
        RECT 661.580 1321.280 661.840 1321.540 ;
        RECT 1807.900 1319.580 1808.160 1319.840 ;
      LAYER met2 ;
        RECT 660.610 1321.650 660.890 1325.025 ;
        RECT 660.610 1321.570 661.780 1321.650 ;
        RECT 660.610 1321.510 661.840 1321.570 ;
        RECT 660.610 1321.025 660.890 1321.510 ;
        RECT 661.580 1321.250 661.840 1321.510 ;
        RECT 1807.900 1319.550 1808.160 1319.870 ;
        RECT 1807.960 17.410 1808.100 1319.550 ;
        RECT 1807.960 17.270 1810.860 17.410 ;
        RECT 1810.720 2.400 1810.860 17.270 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1372.710 32.880 1373.030 32.940 ;
        RECT 1829.030 32.880 1829.350 32.940 ;
        RECT 1372.710 32.740 1829.350 32.880 ;
        RECT 1372.710 32.680 1373.030 32.740 ;
        RECT 1829.030 32.680 1829.350 32.740 ;
      LAYER via ;
        RECT 1372.740 32.680 1373.000 32.940 ;
        RECT 1829.060 32.680 1829.320 32.940 ;
      LAYER met2 ;
        RECT 1370.850 216.650 1371.130 220.000 ;
        RECT 1370.850 216.510 1372.940 216.650 ;
        RECT 1370.850 216.000 1371.130 216.510 ;
        RECT 1372.800 32.970 1372.940 216.510 ;
        RECT 1372.740 32.650 1373.000 32.970 ;
        RECT 1829.060 32.650 1829.320 32.970 ;
        RECT 1829.120 16.050 1829.260 32.650 ;
        RECT 1828.660 15.910 1829.260 16.050 ;
        RECT 1828.660 2.400 1828.800 15.910 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 543.405 1318.265 543.575 1321.495 ;
      LAYER mcon ;
        RECT 543.405 1321.325 543.575 1321.495 ;
      LAYER met1 ;
        RECT 543.330 1321.480 543.650 1321.540 ;
        RECT 543.135 1321.340 543.650 1321.480 ;
        RECT 543.330 1321.280 543.650 1321.340 ;
        RECT 543.345 1318.420 543.635 1318.465 ;
        RECT 1842.370 1318.420 1842.690 1318.480 ;
        RECT 543.345 1318.280 1842.690 1318.420 ;
        RECT 543.345 1318.235 543.635 1318.280 ;
        RECT 1842.370 1318.220 1842.690 1318.280 ;
      LAYER via ;
        RECT 543.360 1321.280 543.620 1321.540 ;
        RECT 1842.400 1318.220 1842.660 1318.480 ;
      LAYER met2 ;
        RECT 541.930 1321.650 542.210 1325.025 ;
        RECT 541.930 1321.570 543.560 1321.650 ;
        RECT 541.930 1321.510 543.620 1321.570 ;
        RECT 541.930 1321.025 542.210 1321.510 ;
        RECT 543.360 1321.250 543.620 1321.510 ;
        RECT 1842.400 1318.190 1842.660 1318.510 ;
        RECT 1842.460 17.410 1842.600 1318.190 ;
        RECT 1842.460 17.270 1846.280 17.410 ;
        RECT 1846.140 2.400 1846.280 17.270 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 710.840 1419.490 710.900 ;
        RECT 1863.070 710.840 1863.390 710.900 ;
        RECT 1419.170 710.700 1863.390 710.840 ;
        RECT 1419.170 710.640 1419.490 710.700 ;
        RECT 1863.070 710.640 1863.390 710.700 ;
      LAYER via ;
        RECT 1419.200 710.640 1419.460 710.900 ;
        RECT 1863.100 710.640 1863.360 710.900 ;
      LAYER met2 ;
        RECT 1419.190 716.875 1419.470 717.245 ;
        RECT 1419.260 710.930 1419.400 716.875 ;
        RECT 1419.200 710.610 1419.460 710.930 ;
        RECT 1863.100 710.610 1863.360 710.930 ;
        RECT 1863.160 17.410 1863.300 710.610 ;
        RECT 1863.160 17.270 1864.220 17.410 ;
        RECT 1864.080 2.400 1864.220 17.270 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
      LAYER via2 ;
        RECT 1419.190 716.920 1419.470 717.200 ;
      LAYER met3 ;
        RECT 1419.165 717.210 1419.495 717.225 ;
        RECT 1408.060 717.120 1419.495 717.210 ;
        RECT 1404.305 716.910 1419.495 717.120 ;
        RECT 1404.305 716.520 1408.305 716.910 ;
        RECT 1419.165 716.895 1419.495 716.910 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 744.810 128.420 745.130 128.480 ;
        RECT 1405.830 128.420 1406.150 128.480 ;
        RECT 744.810 128.280 1406.150 128.420 ;
        RECT 744.810 128.220 745.130 128.280 ;
        RECT 1405.830 128.220 1406.150 128.280 ;
        RECT 740.210 17.240 740.530 17.300 ;
        RECT 744.810 17.240 745.130 17.300 ;
        RECT 740.210 17.100 745.130 17.240 ;
        RECT 740.210 17.040 740.530 17.100 ;
        RECT 744.810 17.040 745.130 17.100 ;
      LAYER via ;
        RECT 744.840 128.220 745.100 128.480 ;
        RECT 1405.860 128.220 1406.120 128.480 ;
        RECT 740.240 17.040 740.500 17.300 ;
        RECT 744.840 17.040 745.100 17.300 ;
      LAYER met2 ;
        RECT 1405.850 421.755 1406.130 422.125 ;
        RECT 1405.920 128.510 1406.060 421.755 ;
        RECT 744.840 128.190 745.100 128.510 ;
        RECT 1405.860 128.190 1406.120 128.510 ;
        RECT 744.900 17.330 745.040 128.190 ;
        RECT 740.240 17.010 740.500 17.330 ;
        RECT 744.840 17.010 745.100 17.330 ;
        RECT 740.300 2.400 740.440 17.010 ;
        RECT 740.090 -4.800 740.650 2.400 ;
      LAYER via2 ;
        RECT 1405.850 421.800 1406.130 422.080 ;
      LAYER met3 ;
        RECT 1404.305 424.120 1408.305 424.720 ;
        RECT 1406.070 422.105 1406.370 424.120 ;
        RECT 1405.825 421.790 1406.370 422.105 ;
        RECT 1405.825 421.775 1406.155 421.790 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 667.605 1319.285 667.775 1321.495 ;
      LAYER mcon ;
        RECT 667.605 1321.325 667.775 1321.495 ;
      LAYER met1 ;
        RECT 667.530 1321.480 667.850 1321.540 ;
        RECT 667.335 1321.340 667.850 1321.480 ;
        RECT 667.530 1321.280 667.850 1321.340 ;
        RECT 667.545 1319.440 667.835 1319.485 ;
        RECT 1876.870 1319.440 1877.190 1319.500 ;
        RECT 667.545 1319.300 1877.190 1319.440 ;
        RECT 667.545 1319.255 667.835 1319.300 ;
        RECT 1876.870 1319.240 1877.190 1319.300 ;
      LAYER via ;
        RECT 667.560 1321.280 667.820 1321.540 ;
        RECT 1876.900 1319.240 1877.160 1319.500 ;
      LAYER met2 ;
        RECT 666.130 1321.650 666.410 1325.025 ;
        RECT 666.130 1321.570 667.760 1321.650 ;
        RECT 666.130 1321.510 667.820 1321.570 ;
        RECT 666.130 1321.025 666.410 1321.510 ;
        RECT 667.560 1321.250 667.820 1321.510 ;
        RECT 1876.900 1319.210 1877.160 1319.530 ;
        RECT 1876.960 17.410 1877.100 1319.210 ;
        RECT 1876.960 17.270 1882.160 17.410 ;
        RECT 1882.020 2.400 1882.160 17.270 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 300.450 182.820 300.770 182.880 ;
        RECT 1897.570 182.820 1897.890 182.880 ;
        RECT 300.450 182.680 1897.890 182.820 ;
        RECT 300.450 182.620 300.770 182.680 ;
        RECT 1897.570 182.620 1897.890 182.680 ;
      LAYER via ;
        RECT 300.480 182.620 300.740 182.880 ;
        RECT 1897.600 182.620 1897.860 182.880 ;
      LAYER met2 ;
        RECT 300.470 395.915 300.750 396.285 ;
        RECT 300.540 182.910 300.680 395.915 ;
        RECT 300.480 182.590 300.740 182.910 ;
        RECT 1897.600 182.590 1897.860 182.910 ;
        RECT 1897.660 17.410 1897.800 182.590 ;
        RECT 1897.660 17.270 1900.100 17.410 ;
        RECT 1899.960 2.400 1900.100 17.270 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
      LAYER via2 ;
        RECT 300.470 395.960 300.750 396.240 ;
      LAYER met3 ;
        RECT 300.445 396.250 300.775 396.265 ;
        RECT 300.445 396.160 310.500 396.250 ;
        RECT 300.445 395.950 314.000 396.160 ;
        RECT 300.445 395.935 300.775 395.950 ;
        RECT 310.000 395.560 314.000 395.950 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 461.910 31.520 462.230 31.580 ;
        RECT 1917.810 31.520 1918.130 31.580 ;
        RECT 461.910 31.380 1918.130 31.520 ;
        RECT 461.910 31.320 462.230 31.380 ;
        RECT 1917.810 31.320 1918.130 31.380 ;
      LAYER via ;
        RECT 461.940 31.320 462.200 31.580 ;
        RECT 1917.840 31.320 1918.100 31.580 ;
      LAYER met2 ;
        RECT 460.970 216.650 461.250 220.000 ;
        RECT 460.970 216.510 462.140 216.650 ;
        RECT 460.970 216.000 461.250 216.510 ;
        RECT 462.000 31.610 462.140 216.510 ;
        RECT 461.940 31.290 462.200 31.610 ;
        RECT 1917.840 31.290 1918.100 31.610 ;
        RECT 1917.900 2.400 1918.040 31.290 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 228.040 1419.490 228.100 ;
        RECT 1932.070 228.040 1932.390 228.100 ;
        RECT 1419.170 227.900 1932.390 228.040 ;
        RECT 1419.170 227.840 1419.490 227.900 ;
        RECT 1932.070 227.840 1932.390 227.900 ;
      LAYER via ;
        RECT 1419.200 227.840 1419.460 228.100 ;
        RECT 1932.100 227.840 1932.360 228.100 ;
      LAYER met2 ;
        RECT 1419.190 234.075 1419.470 234.445 ;
        RECT 1419.260 228.130 1419.400 234.075 ;
        RECT 1419.200 227.810 1419.460 228.130 ;
        RECT 1932.100 227.810 1932.360 228.130 ;
        RECT 1932.160 17.410 1932.300 227.810 ;
        RECT 1932.160 17.270 1935.520 17.410 ;
        RECT 1935.380 2.400 1935.520 17.270 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
      LAYER via2 ;
        RECT 1419.190 234.120 1419.470 234.400 ;
      LAYER met3 ;
        RECT 1419.165 234.410 1419.495 234.425 ;
        RECT 1408.060 234.320 1419.495 234.410 ;
        RECT 1404.305 234.110 1419.495 234.320 ;
        RECT 1404.305 233.720 1408.305 234.110 ;
        RECT 1419.165 234.095 1419.495 234.110 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 672.205 1318.605 672.375 1321.495 ;
      LAYER mcon ;
        RECT 672.205 1321.325 672.375 1321.495 ;
      LAYER met1 ;
        RECT 672.130 1321.480 672.450 1321.540 ;
        RECT 671.935 1321.340 672.450 1321.480 ;
        RECT 672.130 1321.280 672.450 1321.340 ;
        RECT 672.145 1318.760 672.435 1318.805 ;
        RECT 1952.770 1318.760 1953.090 1318.820 ;
        RECT 672.145 1318.620 1953.090 1318.760 ;
        RECT 672.145 1318.575 672.435 1318.620 ;
        RECT 1952.770 1318.560 1953.090 1318.620 ;
      LAYER via ;
        RECT 672.160 1321.280 672.420 1321.540 ;
        RECT 1952.800 1318.560 1953.060 1318.820 ;
      LAYER met2 ;
        RECT 670.730 1321.650 671.010 1325.025 ;
        RECT 670.730 1321.570 672.360 1321.650 ;
        RECT 670.730 1321.510 672.420 1321.570 ;
        RECT 670.730 1321.025 671.010 1321.510 ;
        RECT 672.160 1321.250 672.420 1321.510 ;
        RECT 1952.800 1318.530 1953.060 1318.850 ;
        RECT 1952.860 17.410 1953.000 1318.530 ;
        RECT 1952.860 17.270 1953.460 17.410 ;
        RECT 1953.320 2.400 1953.460 17.270 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1966.570 2.960 1966.890 3.020 ;
        RECT 1971.170 2.960 1971.490 3.020 ;
        RECT 1966.570 2.820 1971.490 2.960 ;
        RECT 1966.570 2.760 1966.890 2.820 ;
        RECT 1971.170 2.760 1971.490 2.820 ;
      LAYER via ;
        RECT 1966.600 2.760 1966.860 3.020 ;
        RECT 1971.200 2.760 1971.460 3.020 ;
      LAYER met2 ;
        RECT 305.530 1243.195 305.810 1243.565 ;
        RECT 305.600 1041.605 305.740 1243.195 ;
        RECT 305.530 1041.235 305.810 1041.605 ;
        RECT 1966.590 106.235 1966.870 106.605 ;
        RECT 1966.660 3.050 1966.800 106.235 ;
        RECT 1966.600 2.730 1966.860 3.050 ;
        RECT 1971.200 2.730 1971.460 3.050 ;
        RECT 1971.260 2.400 1971.400 2.730 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
      LAYER via2 ;
        RECT 305.530 1243.240 305.810 1243.520 ;
        RECT 305.530 1041.280 305.810 1041.560 ;
        RECT 1966.590 106.280 1966.870 106.560 ;
      LAYER met3 ;
        RECT 305.505 1243.530 305.835 1243.545 ;
        RECT 305.505 1243.440 310.500 1243.530 ;
        RECT 305.505 1243.230 314.000 1243.440 ;
        RECT 305.505 1243.215 305.835 1243.230 ;
        RECT 310.000 1242.840 314.000 1243.230 ;
        RECT 305.505 1041.570 305.835 1041.585 ;
        RECT 309.390 1041.570 309.770 1041.580 ;
        RECT 305.505 1041.270 309.770 1041.570 ;
        RECT 305.505 1041.255 305.835 1041.270 ;
        RECT 309.390 1041.260 309.770 1041.270 ;
        RECT 309.390 106.570 309.770 106.580 ;
        RECT 1966.565 106.570 1966.895 106.585 ;
        RECT 309.390 106.270 1966.895 106.570 ;
        RECT 309.390 106.260 309.770 106.270 ;
        RECT 1966.565 106.255 1966.895 106.270 ;
      LAYER via3 ;
        RECT 309.420 1041.260 309.740 1041.580 ;
        RECT 309.420 106.260 309.740 106.580 ;
      LAYER met4 ;
        RECT 309.415 1041.255 309.745 1041.585 ;
        RECT 309.430 106.585 309.730 1041.255 ;
        RECT 309.415 106.255 309.745 106.585 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 273.770 641.820 274.090 641.880 ;
        RECT 296.770 641.820 297.090 641.880 ;
        RECT 273.770 641.680 297.090 641.820 ;
        RECT 273.770 641.620 274.090 641.680 ;
        RECT 296.770 641.620 297.090 641.680 ;
      LAYER via ;
        RECT 273.800 641.620 274.060 641.880 ;
        RECT 296.800 641.620 297.060 641.880 ;
      LAYER met2 ;
        RECT 296.790 643.435 297.070 643.805 ;
        RECT 296.860 641.910 297.000 643.435 ;
        RECT 273.800 641.590 274.060 641.910 ;
        RECT 296.800 641.590 297.060 641.910 ;
        RECT 273.860 45.405 274.000 641.590 ;
        RECT 273.790 45.035 274.070 45.405 ;
        RECT 1989.130 45.035 1989.410 45.405 ;
        RECT 1989.200 2.400 1989.340 45.035 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
      LAYER via2 ;
        RECT 296.790 643.480 297.070 643.760 ;
        RECT 273.790 45.080 274.070 45.360 ;
        RECT 1989.130 45.080 1989.410 45.360 ;
      LAYER met3 ;
        RECT 296.765 643.770 297.095 643.785 ;
        RECT 296.765 643.680 310.500 643.770 ;
        RECT 296.765 643.470 314.000 643.680 ;
        RECT 296.765 643.455 297.095 643.470 ;
        RECT 310.000 643.080 314.000 643.470 ;
        RECT 273.765 45.370 274.095 45.385 ;
        RECT 1989.105 45.370 1989.435 45.385 ;
        RECT 273.765 45.070 1989.435 45.370 ;
        RECT 273.765 45.055 274.095 45.070 ;
        RECT 1989.105 45.055 1989.435 45.070 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 311.030 221.580 311.350 221.640 ;
        RECT 311.030 221.440 1385.360 221.580 ;
        RECT 311.030 221.380 311.350 221.440 ;
        RECT 1385.220 219.600 1385.360 221.440 ;
        RECT 1385.130 219.340 1385.450 219.600 ;
      LAYER via ;
        RECT 311.060 221.380 311.320 221.640 ;
        RECT 1385.160 219.340 1385.420 219.600 ;
      LAYER met2 ;
        RECT 311.050 224.555 311.330 224.925 ;
        RECT 311.120 221.670 311.260 224.555 ;
        RECT 311.060 221.350 311.320 221.670 ;
        RECT 1385.160 219.485 1385.420 219.630 ;
        RECT 1385.150 219.115 1385.430 219.485 ;
        RECT 2006.610 34.155 2006.890 34.525 ;
        RECT 2006.680 2.400 2006.820 34.155 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
      LAYER via2 ;
        RECT 311.050 224.600 311.330 224.880 ;
        RECT 1385.150 219.160 1385.430 219.440 ;
        RECT 2006.610 34.200 2006.890 34.480 ;
      LAYER met3 ;
        RECT 310.000 226.920 314.000 227.520 ;
        RECT 311.270 224.905 311.570 226.920 ;
        RECT 311.025 224.590 311.570 224.905 ;
        RECT 311.025 224.575 311.355 224.590 ;
        RECT 1385.125 219.450 1385.455 219.465 ;
        RECT 1385.790 219.450 1386.170 219.460 ;
        RECT 1385.125 219.150 1386.170 219.450 ;
        RECT 1385.125 219.135 1385.455 219.150 ;
        RECT 1385.790 219.140 1386.170 219.150 ;
        RECT 1385.790 34.490 1386.170 34.500 ;
        RECT 2006.585 34.490 2006.915 34.505 ;
        RECT 1385.790 34.190 2006.915 34.490 ;
        RECT 1385.790 34.180 1386.170 34.190 ;
        RECT 2006.585 34.175 2006.915 34.190 ;
      LAYER via3 ;
        RECT 1385.820 219.140 1386.140 219.460 ;
        RECT 1385.820 34.180 1386.140 34.500 ;
      LAYER met4 ;
        RECT 1385.815 219.135 1386.145 219.465 ;
        RECT 1385.830 34.505 1386.130 219.135 ;
        RECT 1385.815 34.175 1386.145 34.505 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1330.850 33.220 1331.170 33.280 ;
        RECT 2024.530 33.220 2024.850 33.280 ;
        RECT 1330.850 33.080 2024.850 33.220 ;
        RECT 1330.850 33.020 1331.170 33.080 ;
        RECT 2024.530 33.020 2024.850 33.080 ;
      LAYER via ;
        RECT 1330.880 33.020 1331.140 33.280 ;
        RECT 2024.560 33.020 2024.820 33.280 ;
      LAYER met2 ;
        RECT 1331.290 216.650 1331.570 220.000 ;
        RECT 1330.940 216.510 1331.570 216.650 ;
        RECT 1330.940 33.310 1331.080 216.510 ;
        RECT 1331.290 216.000 1331.570 216.510 ;
        RECT 1330.880 32.990 1331.140 33.310 ;
        RECT 2024.560 32.990 2024.820 33.310 ;
        RECT 2024.620 2.400 2024.760 32.990 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1262.310 59.400 1262.630 59.460 ;
        RECT 2042.930 59.400 2043.250 59.460 ;
        RECT 1262.310 59.260 2043.250 59.400 ;
        RECT 1262.310 59.200 1262.630 59.260 ;
        RECT 2042.930 59.200 2043.250 59.260 ;
      LAYER via ;
        RECT 1262.340 59.200 1262.600 59.460 ;
        RECT 2042.960 59.200 2043.220 59.460 ;
      LAYER met2 ;
        RECT 1262.290 216.000 1262.570 220.000 ;
        RECT 1262.400 59.490 1262.540 216.000 ;
        RECT 1262.340 59.170 1262.600 59.490 ;
        RECT 2042.960 59.170 2043.220 59.490 ;
        RECT 2043.020 17.410 2043.160 59.170 ;
        RECT 2042.560 17.270 2043.160 17.410 ;
        RECT 2042.560 2.400 2042.700 17.270 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 753.625 58.225 753.795 137.955 ;
      LAYER mcon ;
        RECT 753.625 137.785 753.795 137.955 ;
      LAYER met1 ;
        RECT 753.090 137.940 753.410 138.000 ;
        RECT 753.565 137.940 753.855 137.985 ;
        RECT 753.090 137.800 753.855 137.940 ;
        RECT 753.090 137.740 753.410 137.800 ;
        RECT 753.565 137.755 753.855 137.800 ;
        RECT 753.550 58.380 753.870 58.440 ;
        RECT 753.355 58.240 753.870 58.380 ;
        RECT 753.550 58.180 753.870 58.240 ;
        RECT 753.550 17.240 753.870 17.300 ;
        RECT 757.690 17.240 758.010 17.300 ;
        RECT 753.550 17.100 758.010 17.240 ;
        RECT 753.550 17.040 753.870 17.100 ;
        RECT 757.690 17.040 758.010 17.100 ;
      LAYER via ;
        RECT 753.120 137.740 753.380 138.000 ;
        RECT 753.580 58.180 753.840 58.440 ;
        RECT 753.580 17.040 753.840 17.300 ;
        RECT 757.720 17.040 757.980 17.300 ;
      LAYER met2 ;
        RECT 757.210 217.330 757.490 220.000 ;
        RECT 755.020 217.190 757.490 217.330 ;
        RECT 755.020 201.690 755.160 217.190 ;
        RECT 757.210 216.000 757.490 217.190 ;
        RECT 754.100 201.550 755.160 201.690 ;
        RECT 754.100 145.365 754.240 201.550 ;
        RECT 753.110 144.995 753.390 145.365 ;
        RECT 754.030 144.995 754.310 145.365 ;
        RECT 753.180 138.030 753.320 144.995 ;
        RECT 753.120 137.710 753.380 138.030 ;
        RECT 753.580 58.150 753.840 58.470 ;
        RECT 753.640 17.330 753.780 58.150 ;
        RECT 753.580 17.010 753.840 17.330 ;
        RECT 757.720 17.010 757.980 17.330 ;
        RECT 757.780 2.400 757.920 17.010 ;
        RECT 757.570 -4.800 758.130 2.400 ;
      LAYER via2 ;
        RECT 753.110 145.040 753.390 145.320 ;
        RECT 754.030 145.040 754.310 145.320 ;
      LAYER met3 ;
        RECT 753.085 145.330 753.415 145.345 ;
        RECT 754.005 145.330 754.335 145.345 ;
        RECT 753.085 145.030 754.335 145.330 ;
        RECT 753.085 145.015 753.415 145.030 ;
        RECT 754.005 145.015 754.335 145.030 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1420.090 538.460 1420.410 538.520 ;
        RECT 2056.270 538.460 2056.590 538.520 ;
        RECT 1420.090 538.320 2056.590 538.460 ;
        RECT 1420.090 538.260 1420.410 538.320 ;
        RECT 2056.270 538.260 2056.590 538.320 ;
      LAYER via ;
        RECT 1420.120 538.260 1420.380 538.520 ;
        RECT 2056.300 538.260 2056.560 538.520 ;
      LAYER met2 ;
        RECT 1420.110 541.435 1420.390 541.805 ;
        RECT 1420.180 538.550 1420.320 541.435 ;
        RECT 1420.120 538.230 1420.380 538.550 ;
        RECT 2056.300 538.230 2056.560 538.550 ;
        RECT 2056.360 16.730 2056.500 538.230 ;
        RECT 2056.360 16.590 2060.640 16.730 ;
        RECT 2060.500 2.400 2060.640 16.590 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
      LAYER via2 ;
        RECT 1420.110 541.480 1420.390 541.760 ;
      LAYER met3 ;
        RECT 1420.085 541.770 1420.415 541.785 ;
        RECT 1408.060 541.680 1420.415 541.770 ;
        RECT 1404.305 541.470 1420.415 541.680 ;
        RECT 1404.305 541.080 1408.305 541.470 ;
        RECT 1420.085 541.455 1420.415 541.470 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2076.970 2.960 2077.290 3.020 ;
        RECT 2078.350 2.960 2078.670 3.020 ;
        RECT 2076.970 2.820 2078.670 2.960 ;
        RECT 2076.970 2.760 2077.290 2.820 ;
        RECT 2078.350 2.760 2078.670 2.820 ;
      LAYER via ;
        RECT 2077.000 2.760 2077.260 3.020 ;
        RECT 2078.380 2.760 2078.640 3.020 ;
      LAYER met2 ;
        RECT 2076.990 168.795 2077.270 169.165 ;
        RECT 2077.060 3.050 2077.200 168.795 ;
        RECT 2077.000 2.730 2077.260 3.050 ;
        RECT 2078.380 2.730 2078.640 3.050 ;
        RECT 2078.440 2.400 2078.580 2.730 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
      LAYER via2 ;
        RECT 2076.990 168.840 2077.270 169.120 ;
      LAYER met3 ;
        RECT 302.950 1053.130 303.330 1053.140 ;
        RECT 302.950 1053.040 310.500 1053.130 ;
        RECT 302.950 1052.830 314.000 1053.040 ;
        RECT 302.950 1052.820 303.330 1052.830 ;
        RECT 310.000 1052.440 314.000 1052.830 ;
        RECT 302.950 169.130 303.330 169.140 ;
        RECT 2076.965 169.130 2077.295 169.145 ;
        RECT 302.950 168.830 2077.295 169.130 ;
        RECT 302.950 168.820 303.330 168.830 ;
        RECT 2076.965 168.815 2077.295 168.830 ;
      LAYER via3 ;
        RECT 302.980 1052.820 303.300 1053.140 ;
        RECT 302.980 168.820 303.300 169.140 ;
      LAYER met4 ;
        RECT 302.975 1052.815 303.305 1053.145 ;
        RECT 302.990 169.145 303.290 1052.815 ;
        RECT 302.975 168.815 303.305 169.145 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 874.070 1347.320 874.390 1347.380 ;
        RECT 2090.770 1347.320 2091.090 1347.380 ;
        RECT 874.070 1347.180 2091.090 1347.320 ;
        RECT 874.070 1347.120 874.390 1347.180 ;
        RECT 2090.770 1347.120 2091.090 1347.180 ;
        RECT 2090.770 2.960 2091.090 3.020 ;
        RECT 2095.830 2.960 2096.150 3.020 ;
        RECT 2090.770 2.820 2096.150 2.960 ;
        RECT 2090.770 2.760 2091.090 2.820 ;
        RECT 2095.830 2.760 2096.150 2.820 ;
      LAYER via ;
        RECT 874.100 1347.120 874.360 1347.380 ;
        RECT 2090.800 1347.120 2091.060 1347.380 ;
        RECT 2090.800 2.760 2091.060 3.020 ;
        RECT 2095.860 2.760 2096.120 3.020 ;
      LAYER met2 ;
        RECT 874.100 1347.090 874.360 1347.410 ;
        RECT 2090.800 1347.090 2091.060 1347.410 ;
        RECT 874.160 1325.025 874.300 1347.090 ;
        RECT 874.050 1321.025 874.330 1325.025 ;
        RECT 2090.860 3.050 2091.000 1347.090 ;
        RECT 2090.800 2.730 2091.060 3.050 ;
        RECT 2095.860 2.730 2096.120 3.050 ;
        RECT 2095.920 2.400 2096.060 2.730 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 663.390 200.500 663.710 200.560 ;
        RECT 668.910 200.500 669.230 200.560 ;
        RECT 663.390 200.360 669.230 200.500 ;
        RECT 663.390 200.300 663.710 200.360 ;
        RECT 668.910 200.300 669.230 200.360 ;
        RECT 668.910 31.860 669.230 31.920 ;
        RECT 2113.770 31.860 2114.090 31.920 ;
        RECT 668.910 31.720 2114.090 31.860 ;
        RECT 668.910 31.660 669.230 31.720 ;
        RECT 2113.770 31.660 2114.090 31.720 ;
      LAYER via ;
        RECT 663.420 200.300 663.680 200.560 ;
        RECT 668.940 200.300 669.200 200.560 ;
        RECT 668.940 31.660 669.200 31.920 ;
        RECT 2113.800 31.660 2114.060 31.920 ;
      LAYER met2 ;
        RECT 663.370 216.000 663.650 220.000 ;
        RECT 663.480 200.590 663.620 216.000 ;
        RECT 663.420 200.270 663.680 200.590 ;
        RECT 668.940 200.270 669.200 200.590 ;
        RECT 669.000 31.950 669.140 200.270 ;
        RECT 668.940 31.630 669.200 31.950 ;
        RECT 2113.800 31.630 2114.060 31.950 ;
        RECT 2113.860 2.400 2114.000 31.630 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 298.150 189.620 298.470 189.680 ;
        RECT 2125.730 189.620 2126.050 189.680 ;
        RECT 298.150 189.480 2126.050 189.620 ;
        RECT 298.150 189.420 298.470 189.480 ;
        RECT 2125.730 189.420 2126.050 189.480 ;
        RECT 2125.730 17.580 2126.050 17.640 ;
        RECT 2131.710 17.580 2132.030 17.640 ;
        RECT 2125.730 17.440 2132.030 17.580 ;
        RECT 2125.730 17.380 2126.050 17.440 ;
        RECT 2131.710 17.380 2132.030 17.440 ;
      LAYER via ;
        RECT 298.180 189.420 298.440 189.680 ;
        RECT 2125.760 189.420 2126.020 189.680 ;
        RECT 2125.760 17.380 2126.020 17.640 ;
        RECT 2131.740 17.380 2132.000 17.640 ;
      LAYER met2 ;
        RECT 298.170 417.675 298.450 418.045 ;
        RECT 298.240 189.710 298.380 417.675 ;
        RECT 298.180 189.390 298.440 189.710 ;
        RECT 2125.760 189.390 2126.020 189.710 ;
        RECT 2125.820 17.670 2125.960 189.390 ;
        RECT 2125.760 17.350 2126.020 17.670 ;
        RECT 2131.740 17.350 2132.000 17.670 ;
        RECT 2131.800 2.400 2131.940 17.350 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
      LAYER via2 ;
        RECT 298.170 417.720 298.450 418.000 ;
      LAYER met3 ;
        RECT 298.145 418.010 298.475 418.025 ;
        RECT 298.145 417.920 310.500 418.010 ;
        RECT 298.145 417.710 314.000 417.920 ;
        RECT 298.145 417.695 298.475 417.710 ;
        RECT 310.000 417.320 314.000 417.710 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 1119.435 306.730 1119.805 ;
        RECT 306.520 966.805 306.660 1119.435 ;
        RECT 306.450 966.435 306.730 966.805 ;
        RECT 2145.990 175.595 2146.270 175.965 ;
        RECT 2146.060 17.410 2146.200 175.595 ;
        RECT 2146.060 17.270 2149.880 17.410 ;
        RECT 2149.740 2.400 2149.880 17.270 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
      LAYER via2 ;
        RECT 306.450 1119.480 306.730 1119.760 ;
        RECT 306.450 966.480 306.730 966.760 ;
        RECT 2145.990 175.640 2146.270 175.920 ;
      LAYER met3 ;
        RECT 306.425 1119.770 306.755 1119.785 ;
        RECT 306.425 1119.680 310.500 1119.770 ;
        RECT 306.425 1119.470 314.000 1119.680 ;
        RECT 306.425 1119.455 306.755 1119.470 ;
        RECT 310.000 1119.080 314.000 1119.470 ;
        RECT 306.425 966.770 306.755 966.785 ;
        RECT 308.470 966.770 308.850 966.780 ;
        RECT 306.425 966.470 308.850 966.770 ;
        RECT 306.425 966.455 306.755 966.470 ;
        RECT 308.470 966.460 308.850 966.470 ;
        RECT 308.470 175.930 308.850 175.940 ;
        RECT 2145.965 175.930 2146.295 175.945 ;
        RECT 308.470 175.630 2146.295 175.930 ;
        RECT 308.470 175.620 308.850 175.630 ;
        RECT 2145.965 175.615 2146.295 175.630 ;
      LAYER via3 ;
        RECT 308.500 966.460 308.820 966.780 ;
        RECT 308.500 175.620 308.820 175.940 ;
      LAYER met4 ;
        RECT 308.495 966.455 308.825 966.785 ;
        RECT 308.510 175.945 308.810 966.455 ;
        RECT 308.495 175.615 308.825 175.945 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 427.960 1419.490 428.020 ;
        RECT 2167.130 427.960 2167.450 428.020 ;
        RECT 1419.170 427.820 2167.450 427.960 ;
        RECT 1419.170 427.760 1419.490 427.820 ;
        RECT 2167.130 427.760 2167.450 427.820 ;
      LAYER via ;
        RECT 1419.200 427.760 1419.460 428.020 ;
        RECT 2167.160 427.760 2167.420 428.020 ;
      LAYER met2 ;
        RECT 1419.190 431.275 1419.470 431.645 ;
        RECT 1419.260 428.050 1419.400 431.275 ;
        RECT 1419.200 427.730 1419.460 428.050 ;
        RECT 2167.160 427.730 2167.420 428.050 ;
        RECT 2167.220 17.410 2167.360 427.730 ;
        RECT 2167.220 17.270 2167.820 17.410 ;
        RECT 2167.680 2.400 2167.820 17.270 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
      LAYER via2 ;
        RECT 1419.190 431.320 1419.470 431.600 ;
      LAYER met3 ;
        RECT 1419.165 431.610 1419.495 431.625 ;
        RECT 1408.060 431.520 1419.495 431.610 ;
        RECT 1404.305 431.310 1419.495 431.520 ;
        RECT 1404.305 430.920 1408.305 431.310 ;
        RECT 1419.165 431.295 1419.495 431.310 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1180.430 1341.200 1180.750 1341.260 ;
        RECT 2180.470 1341.200 2180.790 1341.260 ;
        RECT 1180.430 1341.060 2180.790 1341.200 ;
        RECT 1180.430 1341.000 1180.750 1341.060 ;
        RECT 2180.470 1341.000 2180.790 1341.060 ;
      LAYER via ;
        RECT 1180.460 1341.000 1180.720 1341.260 ;
        RECT 2180.500 1341.000 2180.760 1341.260 ;
      LAYER met2 ;
        RECT 1180.460 1340.970 1180.720 1341.290 ;
        RECT 2180.500 1340.970 2180.760 1341.290 ;
        RECT 1180.520 1325.025 1180.660 1340.970 ;
        RECT 1180.410 1321.025 1180.690 1325.025 ;
        RECT 2180.560 17.410 2180.700 1340.970 ;
        RECT 2180.560 17.270 2185.300 17.410 ;
        RECT 2185.160 2.400 2185.300 17.270 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 599.910 30.840 600.230 30.900 ;
        RECT 2203.010 30.840 2203.330 30.900 ;
        RECT 599.910 30.700 2203.330 30.840 ;
        RECT 599.910 30.640 600.230 30.700 ;
        RECT 2203.010 30.640 2203.330 30.700 ;
      LAYER via ;
        RECT 599.940 30.640 600.200 30.900 ;
        RECT 2203.040 30.640 2203.300 30.900 ;
      LAYER met2 ;
        RECT 598.970 216.650 599.250 220.000 ;
        RECT 598.970 216.510 600.140 216.650 ;
        RECT 598.970 216.000 599.250 216.510 ;
        RECT 600.000 30.930 600.140 216.510 ;
        RECT 599.940 30.610 600.200 30.930 ;
        RECT 2203.040 30.610 2203.300 30.930 ;
        RECT 2203.100 2.400 2203.240 30.610 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 493.190 1353.440 493.510 1353.500 ;
        RECT 2214.970 1353.440 2215.290 1353.500 ;
        RECT 493.190 1353.300 2215.290 1353.440 ;
        RECT 493.190 1353.240 493.510 1353.300 ;
        RECT 2214.970 1353.240 2215.290 1353.300 ;
        RECT 2214.970 16.900 2215.290 16.960 ;
        RECT 2220.950 16.900 2221.270 16.960 ;
        RECT 2214.970 16.760 2221.270 16.900 ;
        RECT 2214.970 16.700 2215.290 16.760 ;
        RECT 2220.950 16.700 2221.270 16.760 ;
      LAYER via ;
        RECT 493.220 1353.240 493.480 1353.500 ;
        RECT 2215.000 1353.240 2215.260 1353.500 ;
        RECT 2215.000 16.700 2215.260 16.960 ;
        RECT 2220.980 16.700 2221.240 16.960 ;
      LAYER met2 ;
        RECT 493.220 1353.210 493.480 1353.530 ;
        RECT 2215.000 1353.210 2215.260 1353.530 ;
        RECT 493.280 1325.025 493.420 1353.210 ;
        RECT 493.170 1321.025 493.450 1325.025 ;
        RECT 2215.060 16.990 2215.200 1353.210 ;
        RECT 2215.000 16.670 2215.260 16.990 ;
        RECT 2220.980 16.670 2221.240 16.990 ;
        RECT 2221.040 2.400 2221.180 16.670 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1313.830 1345.960 1314.150 1346.020 ;
        RECT 1436.190 1345.960 1436.510 1346.020 ;
        RECT 1313.830 1345.820 1436.510 1345.960 ;
        RECT 1313.830 1345.760 1314.150 1345.820 ;
        RECT 1436.190 1345.760 1436.510 1345.820 ;
        RECT 779.310 211.380 779.630 211.440 ;
        RECT 1436.190 211.380 1436.510 211.440 ;
        RECT 779.310 211.240 1436.510 211.380 ;
        RECT 779.310 211.180 779.630 211.240 ;
        RECT 1436.190 211.180 1436.510 211.240 ;
        RECT 775.630 17.240 775.950 17.300 ;
        RECT 779.310 17.240 779.630 17.300 ;
        RECT 775.630 17.100 779.630 17.240 ;
        RECT 775.630 17.040 775.950 17.100 ;
        RECT 779.310 17.040 779.630 17.100 ;
      LAYER via ;
        RECT 1313.860 1345.760 1314.120 1346.020 ;
        RECT 1436.220 1345.760 1436.480 1346.020 ;
        RECT 779.340 211.180 779.600 211.440 ;
        RECT 1436.220 211.180 1436.480 211.440 ;
        RECT 775.660 17.040 775.920 17.300 ;
        RECT 779.340 17.040 779.600 17.300 ;
      LAYER met2 ;
        RECT 1313.860 1345.730 1314.120 1346.050 ;
        RECT 1436.220 1345.730 1436.480 1346.050 ;
        RECT 1313.920 1325.025 1314.060 1345.730 ;
        RECT 1313.810 1321.025 1314.090 1325.025 ;
        RECT 1436.280 211.470 1436.420 1345.730 ;
        RECT 779.340 211.150 779.600 211.470 ;
        RECT 1436.220 211.150 1436.480 211.470 ;
        RECT 779.400 17.330 779.540 211.150 ;
        RECT 775.660 17.010 775.920 17.330 ;
        RECT 779.340 17.010 779.600 17.330 ;
        RECT 775.720 2.400 775.860 17.010 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 855.680 1421.330 855.740 ;
        RECT 2235.670 855.680 2235.990 855.740 ;
        RECT 1421.010 855.540 2235.990 855.680 ;
        RECT 1421.010 855.480 1421.330 855.540 ;
        RECT 2235.670 855.480 2235.990 855.540 ;
      LAYER via ;
        RECT 1421.040 855.480 1421.300 855.740 ;
        RECT 2235.700 855.480 2235.960 855.740 ;
      LAYER met2 ;
        RECT 1421.030 855.595 1421.310 855.965 ;
        RECT 1421.040 855.450 1421.300 855.595 ;
        RECT 2235.700 855.450 2235.960 855.770 ;
        RECT 2235.760 17.410 2235.900 855.450 ;
        RECT 2235.760 17.270 2239.120 17.410 ;
        RECT 2238.980 2.400 2239.120 17.270 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
      LAYER via2 ;
        RECT 1421.030 855.640 1421.310 855.920 ;
      LAYER met3 ;
        RECT 1421.005 855.930 1421.335 855.945 ;
        RECT 1408.060 855.840 1421.335 855.930 ;
        RECT 1404.305 855.630 1421.335 855.840 ;
        RECT 1404.305 855.240 1408.305 855.630 ;
        RECT 1421.005 855.615 1421.335 855.630 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1013.525 1318.945 1013.695 1321.495 ;
      LAYER mcon ;
        RECT 1013.525 1321.325 1013.695 1321.495 ;
      LAYER met1 ;
        RECT 1013.450 1321.480 1013.770 1321.540 ;
        RECT 1013.255 1321.340 1013.770 1321.480 ;
        RECT 1013.450 1321.280 1013.770 1321.340 ;
        RECT 1013.465 1319.100 1013.755 1319.145 ;
        RECT 2256.370 1319.100 2256.690 1319.160 ;
        RECT 1013.465 1318.960 2256.690 1319.100 ;
        RECT 1013.465 1318.915 1013.755 1318.960 ;
        RECT 2256.370 1318.900 2256.690 1318.960 ;
      LAYER via ;
        RECT 1013.480 1321.280 1013.740 1321.540 ;
        RECT 2256.400 1318.900 2256.660 1319.160 ;
      LAYER met2 ;
        RECT 1012.050 1321.650 1012.330 1325.025 ;
        RECT 1012.050 1321.570 1013.680 1321.650 ;
        RECT 1012.050 1321.510 1013.740 1321.570 ;
        RECT 1012.050 1321.025 1012.330 1321.510 ;
        RECT 1013.480 1321.250 1013.740 1321.510 ;
        RECT 2256.400 1318.870 2256.660 1319.190 ;
        RECT 2256.460 2.400 2256.600 1318.870 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 267.330 1083.480 267.650 1083.540 ;
        RECT 297.230 1083.480 297.550 1083.540 ;
        RECT 267.330 1083.340 297.550 1083.480 ;
        RECT 267.330 1083.280 267.650 1083.340 ;
        RECT 297.230 1083.280 297.550 1083.340 ;
      LAYER via ;
        RECT 267.360 1083.280 267.620 1083.540 ;
        RECT 297.260 1083.280 297.520 1083.540 ;
      LAYER met2 ;
        RECT 297.250 1089.515 297.530 1089.885 ;
        RECT 297.320 1083.570 297.460 1089.515 ;
        RECT 267.360 1083.250 267.620 1083.570 ;
        RECT 297.260 1083.250 297.520 1083.570 ;
        RECT 267.420 44.725 267.560 1083.250 ;
        RECT 267.350 44.355 267.630 44.725 ;
        RECT 2274.330 44.355 2274.610 44.725 ;
        RECT 2274.400 2.400 2274.540 44.355 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
      LAYER via2 ;
        RECT 297.250 1089.560 297.530 1089.840 ;
        RECT 267.350 44.400 267.630 44.680 ;
        RECT 2274.330 44.400 2274.610 44.680 ;
      LAYER met3 ;
        RECT 297.225 1089.850 297.555 1089.865 ;
        RECT 297.225 1089.760 310.500 1089.850 ;
        RECT 297.225 1089.550 314.000 1089.760 ;
        RECT 297.225 1089.535 297.555 1089.550 ;
        RECT 310.000 1089.160 314.000 1089.550 ;
        RECT 267.325 44.690 267.655 44.705 ;
        RECT 2274.305 44.690 2274.635 44.705 ;
        RECT 267.325 44.390 2274.635 44.690 ;
        RECT 267.325 44.375 267.655 44.390 ;
        RECT 2274.305 44.375 2274.635 44.390 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 320.230 1353.100 320.550 1353.160 ;
        RECT 2290.870 1353.100 2291.190 1353.160 ;
        RECT 320.230 1352.960 2291.190 1353.100 ;
        RECT 320.230 1352.900 320.550 1352.960 ;
        RECT 2290.870 1352.900 2291.190 1352.960 ;
      LAYER via ;
        RECT 320.260 1352.900 320.520 1353.160 ;
        RECT 2290.900 1352.900 2291.160 1353.160 ;
      LAYER met2 ;
        RECT 320.260 1352.870 320.520 1353.190 ;
        RECT 2290.900 1352.870 2291.160 1353.190 ;
        RECT 320.320 1325.025 320.460 1352.870 ;
        RECT 320.210 1321.025 320.490 1325.025 ;
        RECT 2290.960 17.410 2291.100 1352.870 ;
        RECT 2290.960 17.270 2292.480 17.410 ;
        RECT 2292.340 2.400 2292.480 17.270 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 487.670 1350.040 487.990 1350.100 ;
        RECT 2304.670 1350.040 2304.990 1350.100 ;
        RECT 487.670 1349.900 2304.990 1350.040 ;
        RECT 487.670 1349.840 487.990 1349.900 ;
        RECT 2304.670 1349.840 2304.990 1349.900 ;
      LAYER via ;
        RECT 487.700 1349.840 487.960 1350.100 ;
        RECT 2304.700 1349.840 2304.960 1350.100 ;
      LAYER met2 ;
        RECT 487.700 1349.810 487.960 1350.130 ;
        RECT 2304.700 1349.810 2304.960 1350.130 ;
        RECT 487.760 1325.025 487.900 1349.810 ;
        RECT 487.650 1321.025 487.930 1325.025 ;
        RECT 2304.760 17.410 2304.900 1349.810 ;
        RECT 2304.760 17.270 2310.420 17.410 ;
        RECT 2310.280 2.400 2310.420 17.270 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 819.790 1346.640 820.110 1346.700 ;
        RECT 2325.370 1346.640 2325.690 1346.700 ;
        RECT 819.790 1346.500 2325.690 1346.640 ;
        RECT 819.790 1346.440 820.110 1346.500 ;
        RECT 2325.370 1346.440 2325.690 1346.500 ;
      LAYER via ;
        RECT 819.820 1346.440 820.080 1346.700 ;
        RECT 2325.400 1346.440 2325.660 1346.700 ;
      LAYER met2 ;
        RECT 819.820 1346.410 820.080 1346.730 ;
        RECT 2325.400 1346.410 2325.660 1346.730 ;
        RECT 819.880 1325.025 820.020 1346.410 ;
        RECT 819.770 1321.025 820.050 1325.025 ;
        RECT 2325.460 17.410 2325.600 1346.410 ;
        RECT 2325.460 17.270 2328.360 17.410 ;
        RECT 2328.220 2.400 2328.360 17.270 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 675.350 120.600 675.670 120.660 ;
        RECT 2339.630 120.600 2339.950 120.660 ;
        RECT 675.350 120.460 2339.950 120.600 ;
        RECT 675.350 120.400 675.670 120.460 ;
        RECT 2339.630 120.400 2339.950 120.460 ;
        RECT 2339.630 16.900 2339.950 16.960 ;
        RECT 2345.610 16.900 2345.930 16.960 ;
        RECT 2339.630 16.760 2345.930 16.900 ;
        RECT 2339.630 16.700 2339.950 16.760 ;
        RECT 2345.610 16.700 2345.930 16.760 ;
      LAYER via ;
        RECT 675.380 120.400 675.640 120.660 ;
        RECT 2339.660 120.400 2339.920 120.660 ;
        RECT 2339.660 16.700 2339.920 16.960 ;
        RECT 2345.640 16.700 2345.900 16.960 ;
      LAYER met2 ;
        RECT 673.490 216.650 673.770 220.000 ;
        RECT 673.490 216.510 675.580 216.650 ;
        RECT 673.490 216.000 673.770 216.510 ;
        RECT 675.440 120.690 675.580 216.510 ;
        RECT 675.380 120.370 675.640 120.690 ;
        RECT 2339.660 120.370 2339.920 120.690 ;
        RECT 2339.720 16.990 2339.860 120.370 ;
        RECT 2339.660 16.670 2339.920 16.990 ;
        RECT 2345.640 16.670 2345.900 16.990 ;
        RECT 2345.700 2.400 2345.840 16.670 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2359.890 127.315 2360.170 127.685 ;
        RECT 2359.960 17.410 2360.100 127.315 ;
        RECT 2359.960 17.270 2363.780 17.410 ;
        RECT 2363.640 2.400 2363.780 17.270 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
      LAYER via2 ;
        RECT 2359.890 127.360 2360.170 127.640 ;
      LAYER met3 ;
        RECT 296.510 688.650 296.890 688.660 ;
        RECT 296.510 688.560 310.500 688.650 ;
        RECT 296.510 688.350 314.000 688.560 ;
        RECT 296.510 688.340 296.890 688.350 ;
        RECT 310.000 687.960 314.000 688.350 ;
        RECT 296.510 127.650 296.890 127.660 ;
        RECT 2359.865 127.650 2360.195 127.665 ;
        RECT 296.510 127.350 2360.195 127.650 ;
        RECT 296.510 127.340 296.890 127.350 ;
        RECT 2359.865 127.335 2360.195 127.350 ;
      LAYER via3 ;
        RECT 296.540 688.340 296.860 688.660 ;
        RECT 296.540 127.340 296.860 127.660 ;
      LAYER met4 ;
        RECT 296.535 688.335 296.865 688.665 ;
        RECT 296.550 127.665 296.850 688.335 ;
        RECT 296.535 127.335 296.865 127.665 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 368.990 1352.760 369.310 1352.820 ;
        RECT 2380.570 1352.760 2380.890 1352.820 ;
        RECT 368.990 1352.620 2380.890 1352.760 ;
        RECT 368.990 1352.560 369.310 1352.620 ;
        RECT 2380.570 1352.560 2380.890 1352.620 ;
      LAYER via ;
        RECT 369.020 1352.560 369.280 1352.820 ;
        RECT 2380.600 1352.560 2380.860 1352.820 ;
      LAYER met2 ;
        RECT 369.020 1352.530 369.280 1352.850 ;
        RECT 2380.600 1352.530 2380.860 1352.850 ;
        RECT 369.080 1325.025 369.220 1352.530 ;
        RECT 368.970 1321.025 369.250 1325.025 ;
        RECT 2380.660 17.410 2380.800 1352.530 ;
        RECT 2380.660 17.270 2381.720 17.410 ;
        RECT 2381.580 2.400 2381.720 17.270 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1420.550 1035.200 1420.870 1035.260 ;
        RECT 2394.370 1035.200 2394.690 1035.260 ;
        RECT 1420.550 1035.060 2394.690 1035.200 ;
        RECT 1420.550 1035.000 1420.870 1035.060 ;
        RECT 2394.370 1035.000 2394.690 1035.060 ;
      LAYER via ;
        RECT 1420.580 1035.000 1420.840 1035.260 ;
        RECT 2394.400 1035.000 2394.660 1035.260 ;
      LAYER met2 ;
        RECT 1420.570 1039.195 1420.850 1039.565 ;
        RECT 1420.640 1035.290 1420.780 1039.195 ;
        RECT 1420.580 1034.970 1420.840 1035.290 ;
        RECT 2394.400 1034.970 2394.660 1035.290 ;
        RECT 2394.460 17.410 2394.600 1034.970 ;
        RECT 2394.460 17.270 2399.660 17.410 ;
        RECT 2399.520 2.400 2399.660 17.270 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
      LAYER via2 ;
        RECT 1420.570 1039.240 1420.850 1039.520 ;
      LAYER met3 ;
        RECT 1420.545 1039.530 1420.875 1039.545 ;
        RECT 1408.060 1039.440 1420.875 1039.530 ;
        RECT 1404.305 1039.230 1420.875 1039.440 ;
        RECT 1404.305 1038.840 1408.305 1039.230 ;
        RECT 1420.545 1039.215 1420.875 1039.230 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 793.570 16.900 793.890 16.960 ;
        RECT 800.010 16.900 800.330 16.960 ;
        RECT 793.570 16.760 800.330 16.900 ;
        RECT 793.570 16.700 793.890 16.760 ;
        RECT 800.010 16.700 800.330 16.760 ;
      LAYER via ;
        RECT 793.600 16.700 793.860 16.960 ;
        RECT 800.040 16.700 800.300 16.960 ;
      LAYER met2 ;
        RECT 800.030 79.715 800.310 80.085 ;
        RECT 800.100 16.990 800.240 79.715 ;
        RECT 793.600 16.670 793.860 16.990 ;
        RECT 800.040 16.670 800.300 16.990 ;
        RECT 793.660 2.400 793.800 16.670 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 800.030 79.760 800.310 80.040 ;
      LAYER met3 ;
        RECT 1414.310 1280.250 1414.690 1280.260 ;
        RECT 1408.060 1280.160 1414.690 1280.250 ;
        RECT 1404.305 1279.950 1414.690 1280.160 ;
        RECT 1404.305 1279.560 1408.305 1279.950 ;
        RECT 1414.310 1279.940 1414.690 1279.950 ;
        RECT 800.005 80.050 800.335 80.065 ;
        RECT 1414.310 80.050 1414.690 80.060 ;
        RECT 800.005 79.750 1414.690 80.050 ;
        RECT 800.005 79.735 800.335 79.750 ;
        RECT 1414.310 79.740 1414.690 79.750 ;
      LAYER via3 ;
        RECT 1414.340 1279.940 1414.660 1280.260 ;
        RECT 1414.340 79.740 1414.660 80.060 ;
      LAYER met4 ;
        RECT 1414.335 1279.935 1414.665 1280.265 ;
        RECT 1414.350 80.065 1414.650 1279.935 ;
        RECT 1414.335 79.735 1414.665 80.065 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.310 148.480 641.630 148.540 ;
        RECT 1380.070 148.480 1380.390 148.540 ;
        RECT 641.310 148.340 1380.390 148.480 ;
        RECT 641.310 148.280 641.630 148.340 ;
        RECT 1380.070 148.280 1380.390 148.340 ;
        RECT 639.010 16.560 639.330 16.620 ;
        RECT 641.310 16.560 641.630 16.620 ;
        RECT 639.010 16.420 641.630 16.560 ;
        RECT 639.010 16.360 639.330 16.420 ;
        RECT 641.310 16.360 641.630 16.420 ;
      LAYER via ;
        RECT 641.340 148.280 641.600 148.540 ;
        RECT 1380.100 148.280 1380.360 148.540 ;
        RECT 639.040 16.360 639.300 16.620 ;
        RECT 641.340 16.360 641.600 16.620 ;
      LAYER met2 ;
        RECT 1380.970 216.650 1381.250 220.000 ;
        RECT 1380.160 216.510 1381.250 216.650 ;
        RECT 1380.160 148.570 1380.300 216.510 ;
        RECT 1380.970 216.000 1381.250 216.510 ;
        RECT 641.340 148.250 641.600 148.570 ;
        RECT 1380.100 148.250 1380.360 148.570 ;
        RECT 641.400 16.650 641.540 148.250 ;
        RECT 639.040 16.330 639.300 16.650 ;
        RECT 641.340 16.330 641.600 16.650 ;
        RECT 639.100 2.400 639.240 16.330 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 709.850 141.680 710.170 141.740 ;
        RECT 2421.970 141.680 2422.290 141.740 ;
        RECT 709.850 141.540 2422.290 141.680 ;
        RECT 709.850 141.480 710.170 141.540 ;
        RECT 2421.970 141.480 2422.290 141.540 ;
      LAYER via ;
        RECT 709.880 141.480 710.140 141.740 ;
        RECT 2422.000 141.480 2422.260 141.740 ;
      LAYER met2 ;
        RECT 708.450 216.650 708.730 220.000 ;
        RECT 708.450 216.510 710.080 216.650 ;
        RECT 708.450 216.000 708.730 216.510 ;
        RECT 709.940 141.770 710.080 216.510 ;
        RECT 709.880 141.450 710.140 141.770 ;
        RECT 2422.000 141.450 2422.260 141.770 ;
        RECT 2422.060 17.410 2422.200 141.450 ;
        RECT 2422.060 17.270 2423.120 17.410 ;
        RECT 2422.980 2.400 2423.120 17.270 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 1345.875 374.810 1346.245 ;
        RECT 2435.790 1345.875 2436.070 1346.245 ;
        RECT 374.600 1325.025 374.740 1345.875 ;
        RECT 374.490 1321.025 374.770 1325.025 ;
        RECT 2435.860 17.410 2436.000 1345.875 ;
        RECT 2435.860 17.270 2441.060 17.410 ;
        RECT 2440.920 2.400 2441.060 17.270 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
      LAYER via2 ;
        RECT 374.530 1345.920 374.810 1346.200 ;
        RECT 2435.790 1345.920 2436.070 1346.200 ;
      LAYER met3 ;
        RECT 374.505 1346.210 374.835 1346.225 ;
        RECT 2435.765 1346.210 2436.095 1346.225 ;
        RECT 374.505 1345.910 2436.095 1346.210 ;
        RECT 374.505 1345.895 374.835 1345.910 ;
        RECT 2435.765 1345.895 2436.095 1345.910 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 600.680 1419.490 600.740 ;
        RECT 2456.470 600.680 2456.790 600.740 ;
        RECT 1419.170 600.540 2456.790 600.680 ;
        RECT 1419.170 600.480 1419.490 600.540 ;
        RECT 2456.470 600.480 2456.790 600.540 ;
      LAYER via ;
        RECT 1419.200 600.480 1419.460 600.740 ;
        RECT 2456.500 600.480 2456.760 600.740 ;
      LAYER met2 ;
        RECT 1419.190 606.715 1419.470 607.085 ;
        RECT 1419.260 600.770 1419.400 606.715 ;
        RECT 1419.200 600.450 1419.460 600.770 ;
        RECT 2456.500 600.450 2456.760 600.770 ;
        RECT 2456.560 17.410 2456.700 600.450 ;
        RECT 2456.560 17.270 2459.000 17.410 ;
        RECT 2458.860 2.400 2459.000 17.270 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
      LAYER via2 ;
        RECT 1419.190 606.760 1419.470 607.040 ;
      LAYER met3 ;
        RECT 1419.165 607.050 1419.495 607.065 ;
        RECT 1408.060 606.960 1419.495 607.050 ;
        RECT 1404.305 606.750 1419.495 606.960 ;
        RECT 1404.305 606.360 1408.305 606.750 ;
        RECT 1419.165 606.735 1419.495 606.750 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1131.210 32.200 1131.530 32.260 ;
        RECT 2476.710 32.200 2477.030 32.260 ;
        RECT 1131.210 32.060 2477.030 32.200 ;
        RECT 1131.210 32.000 1131.530 32.060 ;
        RECT 2476.710 32.000 2477.030 32.060 ;
      LAYER via ;
        RECT 1131.240 32.000 1131.500 32.260 ;
        RECT 2476.740 32.000 2477.000 32.260 ;
      LAYER met2 ;
        RECT 1127.970 216.650 1128.250 220.000 ;
        RECT 1127.970 216.510 1131.440 216.650 ;
        RECT 1127.970 216.000 1128.250 216.510 ;
        RECT 1131.300 32.290 1131.440 216.510 ;
        RECT 1131.240 31.970 1131.500 32.290 ;
        RECT 2476.740 31.970 2477.000 32.290 ;
        RECT 2476.800 2.400 2476.940 31.970 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1393.485 1320.305 1393.655 1321.495 ;
      LAYER mcon ;
        RECT 1393.485 1321.325 1393.655 1321.495 ;
      LAYER met1 ;
        RECT 1393.410 1321.480 1393.730 1321.540 ;
        RECT 1393.215 1321.340 1393.730 1321.480 ;
        RECT 1393.410 1321.280 1393.730 1321.340 ;
        RECT 1393.425 1320.460 1393.715 1320.505 ;
        RECT 2490.970 1320.460 2491.290 1320.520 ;
        RECT 1393.425 1320.320 2491.290 1320.460 ;
        RECT 1393.425 1320.275 1393.715 1320.320 ;
        RECT 2490.970 1320.260 2491.290 1320.320 ;
      LAYER via ;
        RECT 1393.440 1321.280 1393.700 1321.540 ;
        RECT 2491.000 1320.260 2491.260 1320.520 ;
      LAYER met2 ;
        RECT 1392.930 1321.650 1393.210 1325.025 ;
        RECT 1392.930 1321.570 1393.640 1321.650 ;
        RECT 1392.930 1321.510 1393.700 1321.570 ;
        RECT 1392.930 1321.025 1393.210 1321.510 ;
        RECT 1393.440 1321.250 1393.700 1321.510 ;
        RECT 2491.000 1320.230 2491.260 1320.550 ;
        RECT 2491.060 17.410 2491.200 1320.230 ;
        RECT 2491.060 17.270 2494.880 17.410 ;
        RECT 2494.740 2.400 2494.880 17.270 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 338.200 1419.490 338.260 ;
        RECT 2480.390 338.200 2480.710 338.260 ;
        RECT 1419.170 338.060 2480.710 338.200 ;
        RECT 1419.170 338.000 1419.490 338.060 ;
        RECT 2480.390 338.000 2480.710 338.060 ;
        RECT 2480.390 17.920 2480.710 17.980 ;
        RECT 2511.670 17.920 2511.990 17.980 ;
        RECT 2480.390 17.780 2511.990 17.920 ;
        RECT 2480.390 17.720 2480.710 17.780 ;
        RECT 2511.670 17.720 2511.990 17.780 ;
      LAYER via ;
        RECT 1419.200 338.000 1419.460 338.260 ;
        RECT 2480.420 338.000 2480.680 338.260 ;
        RECT 2480.420 17.720 2480.680 17.980 ;
        RECT 2511.700 17.720 2511.960 17.980 ;
      LAYER met2 ;
        RECT 1419.190 344.235 1419.470 344.605 ;
        RECT 1419.260 338.290 1419.400 344.235 ;
        RECT 1419.200 337.970 1419.460 338.290 ;
        RECT 2480.420 337.970 2480.680 338.290 ;
        RECT 2480.480 18.010 2480.620 337.970 ;
        RECT 2480.420 17.690 2480.680 18.010 ;
        RECT 2511.700 17.690 2511.960 18.010 ;
        RECT 2511.760 17.410 2511.900 17.690 ;
        RECT 2511.760 17.270 2512.360 17.410 ;
        RECT 2512.220 2.400 2512.360 17.270 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
      LAYER via2 ;
        RECT 1419.190 344.280 1419.470 344.560 ;
      LAYER met3 ;
        RECT 1419.165 344.570 1419.495 344.585 ;
        RECT 1408.060 344.480 1419.495 344.570 ;
        RECT 1404.305 344.270 1419.495 344.480 ;
        RECT 1404.305 343.880 1408.305 344.270 ;
        RECT 1419.165 344.255 1419.495 344.270 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 554.830 200.500 555.150 200.560 ;
        RECT 558.510 200.500 558.830 200.560 ;
        RECT 554.830 200.360 558.830 200.500 ;
        RECT 554.830 200.300 555.150 200.360 ;
        RECT 558.510 200.300 558.830 200.360 ;
        RECT 558.510 86.600 558.830 86.660 ;
        RECT 2525.470 86.600 2525.790 86.660 ;
        RECT 558.510 86.460 2525.790 86.600 ;
        RECT 558.510 86.400 558.830 86.460 ;
        RECT 2525.470 86.400 2525.790 86.460 ;
      LAYER via ;
        RECT 554.860 200.300 555.120 200.560 ;
        RECT 558.540 200.300 558.800 200.560 ;
        RECT 558.540 86.400 558.800 86.660 ;
        RECT 2525.500 86.400 2525.760 86.660 ;
      LAYER met2 ;
        RECT 554.810 216.000 555.090 220.000 ;
        RECT 554.920 200.590 555.060 216.000 ;
        RECT 554.860 200.270 555.120 200.590 ;
        RECT 558.540 200.270 558.800 200.590 ;
        RECT 558.600 86.690 558.740 200.270 ;
        RECT 558.540 86.370 558.800 86.690 ;
        RECT 2525.500 86.370 2525.760 86.690 ;
        RECT 2525.560 17.410 2525.700 86.370 ;
        RECT 2525.560 17.270 2530.300 17.410 ;
        RECT 2530.160 2.400 2530.300 17.270 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1124.960 1421.330 1125.020 ;
        RECT 2487.290 1124.960 2487.610 1125.020 ;
        RECT 1421.010 1124.820 2487.610 1124.960 ;
        RECT 1421.010 1124.760 1421.330 1124.820 ;
        RECT 2487.290 1124.760 2487.610 1124.820 ;
        RECT 2487.290 17.240 2487.610 17.300 ;
        RECT 2548.010 17.240 2548.330 17.300 ;
        RECT 2487.290 17.100 2548.330 17.240 ;
        RECT 2487.290 17.040 2487.610 17.100 ;
        RECT 2548.010 17.040 2548.330 17.100 ;
      LAYER via ;
        RECT 1421.040 1124.760 1421.300 1125.020 ;
        RECT 2487.320 1124.760 2487.580 1125.020 ;
        RECT 2487.320 17.040 2487.580 17.300 ;
        RECT 2548.040 17.040 2548.300 17.300 ;
      LAYER met2 ;
        RECT 1421.030 1126.235 1421.310 1126.605 ;
        RECT 1421.100 1125.050 1421.240 1126.235 ;
        RECT 1421.040 1124.730 1421.300 1125.050 ;
        RECT 2487.320 1124.730 2487.580 1125.050 ;
        RECT 2487.380 17.330 2487.520 1124.730 ;
        RECT 2487.320 17.010 2487.580 17.330 ;
        RECT 2548.040 17.010 2548.300 17.330 ;
        RECT 2548.100 2.400 2548.240 17.010 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1126.280 1421.310 1126.560 ;
      LAYER met3 ;
        RECT 1421.005 1126.570 1421.335 1126.585 ;
        RECT 1408.060 1126.480 1421.335 1126.570 ;
        RECT 1404.305 1126.270 1421.335 1126.480 ;
        RECT 1404.305 1125.880 1408.305 1126.270 ;
        RECT 1421.005 1126.255 1421.335 1126.270 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 1258.155 305.350 1258.525 ;
        RECT 305.140 365.685 305.280 1258.155 ;
        RECT 305.070 365.315 305.350 365.685 ;
        RECT 2560.450 182.395 2560.730 182.765 ;
        RECT 2560.520 17.410 2560.660 182.395 ;
        RECT 2560.520 17.270 2566.180 17.410 ;
        RECT 2566.040 2.400 2566.180 17.270 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
      LAYER via2 ;
        RECT 305.070 1258.200 305.350 1258.480 ;
        RECT 305.070 365.360 305.350 365.640 ;
        RECT 2560.450 182.440 2560.730 182.720 ;
      LAYER met3 ;
        RECT 305.045 1258.490 305.375 1258.505 ;
        RECT 305.045 1258.400 310.500 1258.490 ;
        RECT 305.045 1258.190 314.000 1258.400 ;
        RECT 305.045 1258.175 305.375 1258.190 ;
        RECT 310.000 1257.800 314.000 1258.190 ;
        RECT 305.045 365.650 305.375 365.665 ;
        RECT 307.550 365.650 307.930 365.660 ;
        RECT 305.045 365.350 307.930 365.650 ;
        RECT 305.045 365.335 305.375 365.350 ;
        RECT 307.550 365.340 307.930 365.350 ;
        RECT 307.550 182.730 307.930 182.740 ;
        RECT 2560.425 182.730 2560.755 182.745 ;
        RECT 307.550 182.430 2560.755 182.730 ;
        RECT 307.550 182.420 307.930 182.430 ;
        RECT 2560.425 182.415 2560.755 182.430 ;
      LAYER via3 ;
        RECT 307.580 365.340 307.900 365.660 ;
        RECT 307.580 182.420 307.900 182.740 ;
      LAYER met4 ;
        RECT 307.575 365.335 307.905 365.665 ;
        RECT 307.590 182.745 307.890 365.335 ;
        RECT 307.575 182.415 307.905 182.745 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 890.630 200.500 890.950 200.560 ;
        RECT 896.150 200.500 896.470 200.560 ;
        RECT 890.630 200.360 896.470 200.500 ;
        RECT 890.630 200.300 890.950 200.360 ;
        RECT 896.150 200.300 896.470 200.360 ;
        RECT 896.150 99.860 896.470 99.920 ;
        RECT 2580.670 99.860 2580.990 99.920 ;
        RECT 896.150 99.720 2580.990 99.860 ;
        RECT 896.150 99.660 896.470 99.720 ;
        RECT 2580.670 99.660 2580.990 99.720 ;
      LAYER via ;
        RECT 890.660 200.300 890.920 200.560 ;
        RECT 896.180 200.300 896.440 200.560 ;
        RECT 896.180 99.660 896.440 99.920 ;
        RECT 2580.700 99.660 2580.960 99.920 ;
      LAYER met2 ;
        RECT 890.610 216.000 890.890 220.000 ;
        RECT 890.720 200.590 890.860 216.000 ;
        RECT 890.660 200.270 890.920 200.590 ;
        RECT 896.180 200.270 896.440 200.590 ;
        RECT 896.240 99.950 896.380 200.270 ;
        RECT 896.180 99.630 896.440 99.950 ;
        RECT 2580.700 99.630 2580.960 99.950 ;
        RECT 2580.760 17.410 2580.900 99.630 ;
        RECT 2580.760 17.270 2584.120 17.410 ;
        RECT 2583.980 2.400 2584.120 17.270 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 311.950 175.480 312.270 175.740 ;
        RECT 312.040 174.720 312.180 175.480 ;
        RECT 311.950 174.460 312.270 174.720 ;
        RECT 311.950 99.860 312.270 99.920 ;
        RECT 814.270 99.860 814.590 99.920 ;
        RECT 311.950 99.720 814.590 99.860 ;
        RECT 311.950 99.660 312.270 99.720 ;
        RECT 814.270 99.660 814.590 99.720 ;
      LAYER via ;
        RECT 311.980 175.480 312.240 175.740 ;
        RECT 311.980 174.460 312.240 174.720 ;
        RECT 311.980 99.660 312.240 99.920 ;
        RECT 814.300 99.660 814.560 99.920 ;
      LAYER met2 ;
        RECT 311.970 407.475 312.250 407.845 ;
        RECT 312.040 175.770 312.180 407.475 ;
        RECT 311.980 175.450 312.240 175.770 ;
        RECT 311.980 174.430 312.240 174.750 ;
        RECT 312.040 99.950 312.180 174.430 ;
        RECT 311.980 99.630 312.240 99.950 ;
        RECT 814.300 99.630 814.560 99.950 ;
        RECT 814.360 17.410 814.500 99.630 ;
        RECT 814.360 17.270 817.720 17.410 ;
        RECT 817.580 2.400 817.720 17.270 ;
        RECT 817.370 -4.800 817.930 2.400 ;
      LAYER via2 ;
        RECT 311.970 407.520 312.250 407.800 ;
      LAYER met3 ;
        RECT 310.000 409.160 314.000 409.760 ;
        RECT 312.190 407.825 312.490 409.160 ;
        RECT 311.945 407.510 312.490 407.825 ;
        RECT 311.945 407.495 312.275 407.510 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 906.270 206.280 906.590 206.340 ;
        RECT 910.410 206.280 910.730 206.340 ;
        RECT 906.270 206.140 910.730 206.280 ;
        RECT 906.270 206.080 906.590 206.140 ;
        RECT 910.410 206.080 910.730 206.140 ;
        RECT 910.410 93.740 910.730 93.800 ;
        RECT 2601.830 93.740 2602.150 93.800 ;
        RECT 910.410 93.600 2602.150 93.740 ;
        RECT 910.410 93.540 910.730 93.600 ;
        RECT 2601.830 93.540 2602.150 93.600 ;
      LAYER via ;
        RECT 906.300 206.080 906.560 206.340 ;
        RECT 910.440 206.080 910.700 206.340 ;
        RECT 910.440 93.540 910.700 93.800 ;
        RECT 2601.860 93.540 2602.120 93.800 ;
      LAYER met2 ;
        RECT 906.250 216.000 906.530 220.000 ;
        RECT 906.360 206.370 906.500 216.000 ;
        RECT 906.300 206.050 906.560 206.370 ;
        RECT 910.440 206.050 910.700 206.370 ;
        RECT 910.500 93.830 910.640 206.050 ;
        RECT 910.440 93.510 910.700 93.830 ;
        RECT 2601.860 93.510 2602.120 93.830 ;
        RECT 2601.920 17.410 2602.060 93.510 ;
        RECT 2601.460 17.270 2602.060 17.410 ;
        RECT 2601.460 2.400 2601.600 17.270 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 986.310 24.720 986.630 24.780 ;
        RECT 2619.310 24.720 2619.630 24.780 ;
        RECT 986.310 24.580 2619.630 24.720 ;
        RECT 986.310 24.520 986.630 24.580 ;
        RECT 2619.310 24.520 2619.630 24.580 ;
      LAYER via ;
        RECT 986.340 24.520 986.600 24.780 ;
        RECT 2619.340 24.520 2619.600 24.780 ;
      LAYER met2 ;
        RECT 985.370 216.650 985.650 220.000 ;
        RECT 985.370 216.510 986.540 216.650 ;
        RECT 985.370 216.000 985.650 216.510 ;
        RECT 986.400 24.810 986.540 216.510 ;
        RECT 986.340 24.490 986.600 24.810 ;
        RECT 2619.340 24.490 2619.600 24.810 ;
        RECT 2619.400 2.400 2619.540 24.490 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1295.965 1317.925 1296.135 1322.855 ;
      LAYER mcon ;
        RECT 1295.965 1322.685 1296.135 1322.855 ;
      LAYER met1 ;
        RECT 1295.890 1322.840 1296.210 1322.900 ;
        RECT 1295.695 1322.700 1296.210 1322.840 ;
        RECT 1295.890 1322.640 1296.210 1322.700 ;
        RECT 1295.905 1318.080 1296.195 1318.125 ;
        RECT 2635.870 1318.080 2636.190 1318.140 ;
        RECT 1295.905 1317.940 2636.190 1318.080 ;
        RECT 1295.905 1317.895 1296.195 1317.940 ;
        RECT 2635.870 1317.880 2636.190 1317.940 ;
      LAYER via ;
        RECT 1295.920 1322.640 1296.180 1322.900 ;
        RECT 2635.900 1317.880 2636.160 1318.140 ;
      LAYER met2 ;
        RECT 1294.490 1323.010 1294.770 1325.025 ;
        RECT 1294.490 1322.930 1296.120 1323.010 ;
        RECT 1294.490 1322.870 1296.180 1322.930 ;
        RECT 1294.490 1321.025 1294.770 1322.870 ;
        RECT 1295.920 1322.610 1296.180 1322.870 ;
        RECT 2635.900 1317.850 2636.160 1318.170 ;
        RECT 2635.960 17.410 2636.100 1317.850 ;
        RECT 2635.960 17.270 2637.480 17.410 ;
        RECT 2637.340 2.400 2637.480 17.270 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 1184.715 302.590 1185.085 ;
        RECT 302.380 379.285 302.520 1184.715 ;
        RECT 302.310 378.915 302.590 379.285 ;
        RECT 2649.690 162.675 2649.970 163.045 ;
        RECT 2649.760 17.410 2649.900 162.675 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
      LAYER via2 ;
        RECT 302.310 1184.760 302.590 1185.040 ;
        RECT 302.310 378.960 302.590 379.240 ;
        RECT 2649.690 162.720 2649.970 163.000 ;
      LAYER met3 ;
        RECT 302.285 1185.050 302.615 1185.065 ;
        RECT 302.285 1184.960 310.500 1185.050 ;
        RECT 302.285 1184.750 314.000 1184.960 ;
        RECT 302.285 1184.735 302.615 1184.750 ;
        RECT 310.000 1184.360 314.000 1184.750 ;
        RECT 302.285 379.260 302.615 379.265 ;
        RECT 302.030 379.250 302.615 379.260 ;
        RECT 301.830 378.950 302.615 379.250 ;
        RECT 302.030 378.940 302.615 378.950 ;
        RECT 302.285 378.935 302.615 378.940 ;
        RECT 302.030 163.010 302.410 163.020 ;
        RECT 2649.665 163.010 2649.995 163.025 ;
        RECT 302.030 162.710 2649.995 163.010 ;
        RECT 302.030 162.700 302.410 162.710 ;
        RECT 2649.665 162.695 2649.995 162.710 ;
      LAYER via3 ;
        RECT 302.060 378.940 302.380 379.260 ;
        RECT 302.060 162.700 302.380 163.020 ;
      LAYER met4 ;
        RECT 302.055 378.935 302.385 379.265 ;
        RECT 302.070 163.025 302.370 378.935 ;
        RECT 302.055 162.695 302.385 163.025 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 358.940 1421.330 359.000 ;
        RECT 1673.090 358.940 1673.410 359.000 ;
        RECT 1421.010 358.800 1673.410 358.940 ;
        RECT 1421.010 358.740 1421.330 358.800 ;
        RECT 1673.090 358.740 1673.410 358.800 ;
        RECT 1673.090 217.500 1673.410 217.560 ;
        RECT 2670.370 217.500 2670.690 217.560 ;
        RECT 1673.090 217.360 2670.690 217.500 ;
        RECT 1673.090 217.300 1673.410 217.360 ;
        RECT 2670.370 217.300 2670.690 217.360 ;
      LAYER via ;
        RECT 1421.040 358.740 1421.300 359.000 ;
        RECT 1673.120 358.740 1673.380 359.000 ;
        RECT 1673.120 217.300 1673.380 217.560 ;
        RECT 2670.400 217.300 2670.660 217.560 ;
      LAYER met2 ;
        RECT 1421.030 359.195 1421.310 359.565 ;
        RECT 1421.100 359.030 1421.240 359.195 ;
        RECT 1421.040 358.710 1421.300 359.030 ;
        RECT 1673.120 358.710 1673.380 359.030 ;
        RECT 1673.180 217.590 1673.320 358.710 ;
        RECT 1673.120 217.270 1673.380 217.590 ;
        RECT 2670.400 217.270 2670.660 217.590 ;
        RECT 2670.460 17.410 2670.600 217.270 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
      LAYER via2 ;
        RECT 1421.030 359.240 1421.310 359.520 ;
      LAYER met3 ;
        RECT 1421.005 359.530 1421.335 359.545 ;
        RECT 1408.060 359.440 1421.335 359.530 ;
        RECT 1404.305 359.230 1421.335 359.440 ;
        RECT 1404.305 358.840 1408.305 359.230 ;
        RECT 1421.005 359.215 1421.335 359.230 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1069.110 38.660 1069.430 38.720 ;
        RECT 2690.610 38.660 2690.930 38.720 ;
        RECT 1069.110 38.520 2690.930 38.660 ;
        RECT 1069.110 38.460 1069.430 38.520 ;
        RECT 2690.610 38.460 2690.930 38.520 ;
      LAYER via ;
        RECT 1069.140 38.460 1069.400 38.720 ;
        RECT 2690.640 38.460 2690.900 38.720 ;
      LAYER met2 ;
        RECT 1069.090 216.000 1069.370 220.000 ;
        RECT 1069.200 38.750 1069.340 216.000 ;
        RECT 1069.140 38.430 1069.400 38.750 ;
        RECT 2690.640 38.430 2690.900 38.750 ;
        RECT 2690.700 2.400 2690.840 38.430 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1206.650 31.180 1206.970 31.240 ;
        RECT 2708.550 31.180 2708.870 31.240 ;
        RECT 1206.650 31.040 2708.870 31.180 ;
        RECT 1206.650 30.980 1206.970 31.040 ;
        RECT 2708.550 30.980 2708.870 31.040 ;
      LAYER via ;
        RECT 1206.680 30.980 1206.940 31.240 ;
        RECT 2708.580 30.980 2708.840 31.240 ;
      LAYER met2 ;
        RECT 1207.090 216.650 1207.370 220.000 ;
        RECT 1206.740 216.510 1207.370 216.650 ;
        RECT 1206.740 31.270 1206.880 216.510 ;
        RECT 1207.090 216.000 1207.370 216.510 ;
        RECT 1206.680 30.950 1206.940 31.270 ;
        RECT 2708.580 30.950 2708.840 31.270 ;
        RECT 2708.640 2.400 2708.780 30.950 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1124.310 39.000 1124.630 39.060 ;
        RECT 2726.490 39.000 2726.810 39.060 ;
        RECT 1124.310 38.860 2726.810 39.000 ;
        RECT 1124.310 38.800 1124.630 38.860 ;
        RECT 2726.490 38.800 2726.810 38.860 ;
      LAYER via ;
        RECT 1124.340 38.800 1124.600 39.060 ;
        RECT 2726.520 38.800 2726.780 39.060 ;
      LAYER met2 ;
        RECT 1123.370 216.650 1123.650 220.000 ;
        RECT 1123.370 216.510 1124.540 216.650 ;
        RECT 1123.370 216.000 1123.650 216.510 ;
        RECT 1124.400 39.090 1124.540 216.510 ;
        RECT 1124.340 38.770 1124.600 39.090 ;
        RECT 2726.520 38.770 2726.780 39.090 ;
        RECT 2726.580 2.400 2726.720 38.770 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1165.250 1325.220 1165.570 1325.280 ;
        RECT 2739.370 1325.220 2739.690 1325.280 ;
        RECT 1165.250 1325.080 2739.690 1325.220 ;
        RECT 1165.250 1325.020 1165.570 1325.080 ;
        RECT 2739.370 1325.020 2739.690 1325.080 ;
        RECT 2739.370 2.960 2739.690 3.020 ;
        RECT 2744.430 2.960 2744.750 3.020 ;
        RECT 2739.370 2.820 2744.750 2.960 ;
        RECT 2739.370 2.760 2739.690 2.820 ;
        RECT 2744.430 2.760 2744.750 2.820 ;
      LAYER via ;
        RECT 1165.280 1325.020 1165.540 1325.280 ;
        RECT 2739.400 1325.020 2739.660 1325.280 ;
        RECT 2739.400 2.760 2739.660 3.020 ;
        RECT 2744.460 2.760 2744.720 3.020 ;
      LAYER met2 ;
        RECT 1165.280 1325.050 1165.540 1325.310 ;
        RECT 1165.280 1325.025 1165.870 1325.050 ;
        RECT 1165.280 1324.990 1165.970 1325.025 ;
        RECT 2739.400 1324.990 2739.660 1325.310 ;
        RECT 1165.340 1324.910 1165.970 1324.990 ;
        RECT 1165.690 1321.025 1165.970 1324.910 ;
        RECT 2739.460 3.050 2739.600 1324.990 ;
        RECT 2739.400 2.730 2739.660 3.050 ;
        RECT 2744.460 2.730 2744.720 3.050 ;
        RECT 2744.520 2.400 2744.660 2.730 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 883.560 1421.330 883.620 ;
        RECT 2514.890 883.560 2515.210 883.620 ;
        RECT 1421.010 883.420 2515.210 883.560 ;
        RECT 1421.010 883.360 1421.330 883.420 ;
        RECT 2514.890 883.360 2515.210 883.420 ;
        RECT 2514.890 18.600 2515.210 18.660 ;
        RECT 2514.890 18.460 2518.800 18.600 ;
        RECT 2514.890 18.400 2515.210 18.460 ;
        RECT 2518.660 17.920 2518.800 18.460 ;
        RECT 2761.910 17.920 2762.230 17.980 ;
        RECT 2518.660 17.780 2762.230 17.920 ;
        RECT 2761.910 17.720 2762.230 17.780 ;
      LAYER via ;
        RECT 1421.040 883.360 1421.300 883.620 ;
        RECT 2514.920 883.360 2515.180 883.620 ;
        RECT 2514.920 18.400 2515.180 18.660 ;
        RECT 2761.940 17.720 2762.200 17.980 ;
      LAYER met2 ;
        RECT 1421.030 885.515 1421.310 885.885 ;
        RECT 1421.100 883.650 1421.240 885.515 ;
        RECT 1421.040 883.330 1421.300 883.650 ;
        RECT 2514.920 883.330 2515.180 883.650 ;
        RECT 2514.980 18.690 2515.120 883.330 ;
        RECT 2514.920 18.370 2515.180 18.690 ;
        RECT 2761.940 17.690 2762.200 18.010 ;
        RECT 2762.000 2.400 2762.140 17.690 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
      LAYER via2 ;
        RECT 1421.030 885.560 1421.310 885.840 ;
      LAYER met3 ;
        RECT 1421.005 885.850 1421.335 885.865 ;
        RECT 1408.060 885.760 1421.335 885.850 ;
        RECT 1404.305 885.550 1421.335 885.760 ;
        RECT 1404.305 885.160 1408.305 885.550 ;
        RECT 1421.005 885.535 1421.335 885.550 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 678.110 200.500 678.430 200.560 ;
        RECT 682.250 200.500 682.570 200.560 ;
        RECT 678.110 200.360 682.570 200.500 ;
        RECT 678.110 200.300 678.430 200.360 ;
        RECT 682.250 200.300 682.570 200.360 ;
        RECT 682.250 60.080 682.570 60.140 ;
        RECT 834.970 60.080 835.290 60.140 ;
        RECT 682.250 59.940 835.290 60.080 ;
        RECT 682.250 59.880 682.570 59.940 ;
        RECT 834.970 59.880 835.290 59.940 ;
      LAYER via ;
        RECT 678.140 200.300 678.400 200.560 ;
        RECT 682.280 200.300 682.540 200.560 ;
        RECT 682.280 59.880 682.540 60.140 ;
        RECT 835.000 59.880 835.260 60.140 ;
      LAYER met2 ;
        RECT 678.090 216.000 678.370 220.000 ;
        RECT 678.200 200.590 678.340 216.000 ;
        RECT 678.140 200.270 678.400 200.590 ;
        RECT 682.280 200.270 682.540 200.590 ;
        RECT 682.340 60.170 682.480 200.270 ;
        RECT 682.280 59.850 682.540 60.170 ;
        RECT 835.000 59.850 835.260 60.170 ;
        RECT 835.060 17.410 835.200 59.850 ;
        RECT 835.060 17.270 835.660 17.410 ;
        RECT 835.520 2.400 835.660 17.270 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1020.810 37.980 1021.130 38.040 ;
        RECT 2779.850 37.980 2780.170 38.040 ;
        RECT 1020.810 37.840 2780.170 37.980 ;
        RECT 1020.810 37.780 1021.130 37.840 ;
        RECT 2779.850 37.780 2780.170 37.840 ;
      LAYER via ;
        RECT 1020.840 37.780 1021.100 38.040 ;
        RECT 2779.880 37.780 2780.140 38.040 ;
      LAYER met2 ;
        RECT 1019.410 216.650 1019.690 220.000 ;
        RECT 1019.410 216.510 1021.040 216.650 ;
        RECT 1019.410 216.000 1019.690 216.510 ;
        RECT 1020.900 38.070 1021.040 216.510 ;
        RECT 1020.840 37.750 1021.100 38.070 ;
        RECT 2779.880 37.750 2780.140 38.070 ;
        RECT 2779.940 2.400 2780.080 37.750 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 346.910 200.500 347.230 200.560 ;
        RECT 351.510 200.500 351.830 200.560 ;
        RECT 346.910 200.360 351.830 200.500 ;
        RECT 346.910 200.300 347.230 200.360 ;
        RECT 351.510 200.300 351.830 200.360 ;
        RECT 351.510 134.540 351.830 134.600 ;
        RECT 2794.570 134.540 2794.890 134.600 ;
        RECT 351.510 134.400 2794.890 134.540 ;
        RECT 351.510 134.340 351.830 134.400 ;
        RECT 2794.570 134.340 2794.890 134.400 ;
      LAYER via ;
        RECT 346.940 200.300 347.200 200.560 ;
        RECT 351.540 200.300 351.800 200.560 ;
        RECT 351.540 134.340 351.800 134.600 ;
        RECT 2794.600 134.340 2794.860 134.600 ;
      LAYER met2 ;
        RECT 346.890 216.000 347.170 220.000 ;
        RECT 347.000 200.590 347.140 216.000 ;
        RECT 346.940 200.270 347.200 200.590 ;
        RECT 351.540 200.270 351.800 200.590 ;
        RECT 351.600 134.630 351.740 200.270 ;
        RECT 351.540 134.310 351.800 134.630 ;
        RECT 2794.600 134.310 2794.860 134.630 ;
        RECT 2794.660 17.410 2794.800 134.310 ;
        RECT 2794.660 17.270 2798.020 17.410 ;
        RECT 2797.880 2.400 2798.020 17.270 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1344.650 148.140 1344.970 148.200 ;
        RECT 2815.270 148.140 2815.590 148.200 ;
        RECT 1344.650 148.000 2815.590 148.140 ;
        RECT 1344.650 147.940 1344.970 148.000 ;
        RECT 2815.270 147.940 2815.590 148.000 ;
      LAYER via ;
        RECT 1344.680 147.940 1344.940 148.200 ;
        RECT 2815.300 147.940 2815.560 148.200 ;
      LAYER met2 ;
        RECT 1341.410 216.650 1341.690 220.000 ;
        RECT 1341.410 216.510 1344.880 216.650 ;
        RECT 1341.410 216.000 1341.690 216.510 ;
        RECT 1344.740 148.230 1344.880 216.510 ;
        RECT 1344.680 147.910 1344.940 148.230 ;
        RECT 2815.300 147.910 2815.560 148.230 ;
        RECT 2815.360 17.410 2815.500 147.910 ;
        RECT 2815.360 17.270 2815.960 17.410 ;
        RECT 2815.820 2.400 2815.960 17.270 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 339.550 1333.380 339.870 1333.440 ;
        RECT 634.870 1333.380 635.190 1333.440 ;
        RECT 339.550 1333.240 635.190 1333.380 ;
        RECT 339.550 1333.180 339.870 1333.240 ;
        RECT 634.870 1333.180 635.190 1333.240 ;
      LAYER via ;
        RECT 339.580 1333.180 339.840 1333.440 ;
        RECT 634.900 1333.180 635.160 1333.440 ;
      LAYER met2 ;
        RECT 339.580 1333.150 339.840 1333.470 ;
        RECT 634.900 1333.150 635.160 1333.470 ;
        RECT 339.640 1325.025 339.780 1333.150 ;
        RECT 634.960 1327.885 635.100 1333.150 ;
        RECT 634.890 1327.515 635.170 1327.885 ;
        RECT 2829.090 1327.515 2829.370 1327.885 ;
        RECT 339.530 1321.025 339.810 1325.025 ;
        RECT 2829.160 17.410 2829.300 1327.515 ;
        RECT 2829.160 17.270 2833.900 17.410 ;
        RECT 2833.760 2.400 2833.900 17.270 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
      LAYER via2 ;
        RECT 634.890 1327.560 635.170 1327.840 ;
        RECT 2829.090 1327.560 2829.370 1327.840 ;
      LAYER met3 ;
        RECT 634.865 1327.850 635.195 1327.865 ;
        RECT 2829.065 1327.850 2829.395 1327.865 ;
        RECT 634.865 1327.550 2829.395 1327.850 ;
        RECT 634.865 1327.535 635.195 1327.550 ;
        RECT 2829.065 1327.535 2829.395 1327.550 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 606.810 72.320 607.130 72.380 ;
        RECT 2849.770 72.320 2850.090 72.380 ;
        RECT 606.810 72.180 2850.090 72.320 ;
        RECT 606.810 72.120 607.130 72.180 ;
        RECT 2849.770 72.120 2850.090 72.180 ;
      LAYER via ;
        RECT 606.840 72.120 607.100 72.380 ;
        RECT 2849.800 72.120 2850.060 72.380 ;
      LAYER met2 ;
        RECT 604.490 216.650 604.770 220.000 ;
        RECT 604.490 216.510 607.040 216.650 ;
        RECT 604.490 216.000 604.770 216.510 ;
        RECT 606.900 72.410 607.040 216.510 ;
        RECT 606.840 72.090 607.100 72.410 ;
        RECT 2849.800 72.090 2850.060 72.410 ;
        RECT 2849.860 17.410 2850.000 72.090 ;
        RECT 2849.860 17.270 2851.380 17.410 ;
        RECT 2851.240 2.400 2851.380 17.270 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 856.590 200.500 856.910 200.560 ;
        RECT 861.650 200.500 861.970 200.560 ;
        RECT 856.590 200.360 861.970 200.500 ;
        RECT 856.590 200.300 856.910 200.360 ;
        RECT 861.650 200.300 861.970 200.360 ;
        RECT 861.650 168.880 861.970 168.940 ;
        RECT 2863.570 168.880 2863.890 168.940 ;
        RECT 861.650 168.740 2863.890 168.880 ;
        RECT 861.650 168.680 861.970 168.740 ;
        RECT 2863.570 168.680 2863.890 168.740 ;
      LAYER via ;
        RECT 856.620 200.300 856.880 200.560 ;
        RECT 861.680 200.300 861.940 200.560 ;
        RECT 861.680 168.680 861.940 168.940 ;
        RECT 2863.600 168.680 2863.860 168.940 ;
      LAYER met2 ;
        RECT 856.570 216.000 856.850 220.000 ;
        RECT 856.680 200.590 856.820 216.000 ;
        RECT 856.620 200.270 856.880 200.590 ;
        RECT 861.680 200.270 861.940 200.590 ;
        RECT 861.740 168.970 861.880 200.270 ;
        RECT 861.680 168.650 861.940 168.970 ;
        RECT 2863.600 168.650 2863.860 168.970 ;
        RECT 2863.660 17.410 2863.800 168.650 ;
        RECT 2863.660 17.270 2869.320 17.410 ;
        RECT 2869.180 2.400 2869.320 17.270 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1076.680 1421.330 1076.740 ;
        RECT 2570.090 1076.680 2570.410 1076.740 ;
        RECT 1421.010 1076.540 2570.410 1076.680 ;
        RECT 1421.010 1076.480 1421.330 1076.540 ;
        RECT 2570.090 1076.480 2570.410 1076.540 ;
        RECT 2570.090 20.640 2570.410 20.700 ;
        RECT 2572.850 20.640 2573.170 20.700 ;
        RECT 2570.090 20.500 2573.170 20.640 ;
        RECT 2570.090 20.440 2570.410 20.500 ;
        RECT 2572.850 20.440 2573.170 20.500 ;
        RECT 2572.850 17.240 2573.170 17.300 ;
        RECT 2887.030 17.240 2887.350 17.300 ;
        RECT 2572.850 17.100 2887.350 17.240 ;
        RECT 2572.850 17.040 2573.170 17.100 ;
        RECT 2887.030 17.040 2887.350 17.100 ;
      LAYER via ;
        RECT 1421.040 1076.480 1421.300 1076.740 ;
        RECT 2570.120 1076.480 2570.380 1076.740 ;
        RECT 2570.120 20.440 2570.380 20.700 ;
        RECT 2572.880 20.440 2573.140 20.700 ;
        RECT 2572.880 17.040 2573.140 17.300 ;
        RECT 2887.060 17.040 2887.320 17.300 ;
      LAYER met2 ;
        RECT 1421.030 1082.715 1421.310 1083.085 ;
        RECT 1421.100 1076.770 1421.240 1082.715 ;
        RECT 1421.040 1076.450 1421.300 1076.770 ;
        RECT 2570.120 1076.450 2570.380 1076.770 ;
        RECT 2570.180 20.730 2570.320 1076.450 ;
        RECT 2570.120 20.410 2570.380 20.730 ;
        RECT 2572.880 20.410 2573.140 20.730 ;
        RECT 2572.940 17.330 2573.080 20.410 ;
        RECT 2572.880 17.010 2573.140 17.330 ;
        RECT 2887.060 17.010 2887.320 17.330 ;
        RECT 2887.120 2.400 2887.260 17.010 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1082.760 1421.310 1083.040 ;
      LAYER met3 ;
        RECT 1421.005 1083.050 1421.335 1083.065 ;
        RECT 1408.060 1082.960 1421.335 1083.050 ;
        RECT 1404.305 1082.750 1421.335 1082.960 ;
        RECT 1404.305 1082.360 1408.305 1082.750 ;
        RECT 1421.005 1082.735 1421.335 1082.750 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2873.690 17.580 2874.010 17.640 ;
        RECT 2904.970 17.580 2905.290 17.640 ;
        RECT 2873.690 17.440 2905.290 17.580 ;
        RECT 2873.690 17.380 2874.010 17.440 ;
        RECT 2904.970 17.380 2905.290 17.440 ;
      LAYER via ;
        RECT 2873.720 17.380 2873.980 17.640 ;
        RECT 2905.000 17.380 2905.260 17.640 ;
      LAYER met2 ;
        RECT 572.330 1325.475 572.610 1325.845 ;
        RECT 2873.710 1325.475 2873.990 1325.845 ;
        RECT 572.400 1325.025 572.540 1325.475 ;
        RECT 572.290 1321.025 572.570 1325.025 ;
        RECT 2873.780 17.670 2873.920 1325.475 ;
        RECT 2873.720 17.350 2873.980 17.670 ;
        RECT 2905.000 17.350 2905.260 17.670 ;
        RECT 2905.060 2.400 2905.200 17.350 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 572.330 1325.520 572.610 1325.800 ;
        RECT 2873.710 1325.520 2873.990 1325.800 ;
      LAYER met3 ;
        RECT 572.305 1325.810 572.635 1325.825 ;
        RECT 2873.685 1325.810 2874.015 1325.825 ;
        RECT 572.305 1325.510 2874.015 1325.810 ;
        RECT 572.305 1325.495 572.635 1325.510 ;
        RECT 2873.685 1325.495 2874.015 1325.510 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 854.750 128.760 855.070 128.820 ;
        RECT 1410.430 128.760 1410.750 128.820 ;
        RECT 854.750 128.620 1410.750 128.760 ;
        RECT 854.750 128.560 855.070 128.620 ;
        RECT 1410.430 128.560 1410.750 128.620 ;
      LAYER via ;
        RECT 854.780 128.560 855.040 128.820 ;
        RECT 1410.460 128.560 1410.720 128.820 ;
      LAYER met2 ;
        RECT 1410.450 380.955 1410.730 381.325 ;
        RECT 1410.520 128.850 1410.660 380.955 ;
        RECT 854.780 128.530 855.040 128.850 ;
        RECT 1410.460 128.530 1410.720 128.850 ;
        RECT 854.840 17.410 854.980 128.530 ;
        RECT 853.000 17.270 854.980 17.410 ;
        RECT 853.000 2.400 853.140 17.270 ;
        RECT 852.790 -4.800 853.350 2.400 ;
      LAYER via2 ;
        RECT 1410.450 381.000 1410.730 381.280 ;
      LAYER met3 ;
        RECT 1410.425 381.290 1410.755 381.305 ;
        RECT 1408.060 381.200 1410.755 381.290 ;
        RECT 1404.305 380.990 1410.755 381.200 ;
        RECT 1404.305 380.600 1408.305 380.990 ;
        RECT 1410.425 380.975 1410.755 380.990 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.690 216.650 866.970 220.000 ;
        RECT 866.690 216.510 869.240 216.650 ;
        RECT 866.690 216.000 866.970 216.510 ;
        RECT 869.100 103.090 869.240 216.510 ;
        RECT 869.100 102.950 869.700 103.090 ;
        RECT 869.560 17.410 869.700 102.950 ;
        RECT 869.560 17.270 871.080 17.410 ;
        RECT 870.940 2.400 871.080 17.270 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 738.445 1317.925 738.615 1321.495 ;
      LAYER mcon ;
        RECT 738.445 1321.325 738.615 1321.495 ;
      LAYER met1 ;
        RECT 738.370 1321.480 738.690 1321.540 ;
        RECT 738.175 1321.340 738.690 1321.480 ;
        RECT 738.370 1321.280 738.690 1321.340 ;
        RECT 268.250 1318.080 268.570 1318.140 ;
        RECT 738.385 1318.080 738.675 1318.125 ;
        RECT 268.250 1317.940 738.675 1318.080 ;
        RECT 268.250 1317.880 268.570 1317.940 ;
        RECT 738.385 1317.895 738.675 1317.940 ;
        RECT 268.250 33.220 268.570 33.280 ;
        RECT 888.790 33.220 889.110 33.280 ;
        RECT 268.250 33.080 889.110 33.220 ;
        RECT 268.250 33.020 268.570 33.080 ;
        RECT 888.790 33.020 889.110 33.080 ;
      LAYER via ;
        RECT 738.400 1321.280 738.660 1321.540 ;
        RECT 268.280 1317.880 268.540 1318.140 ;
        RECT 268.280 33.020 268.540 33.280 ;
        RECT 888.820 33.020 889.080 33.280 ;
      LAYER met2 ;
        RECT 739.730 1321.650 740.010 1325.025 ;
        RECT 738.460 1321.570 740.010 1321.650 ;
        RECT 738.400 1321.510 740.010 1321.570 ;
        RECT 738.400 1321.250 738.660 1321.510 ;
        RECT 739.730 1321.025 740.010 1321.510 ;
        RECT 268.280 1317.850 268.540 1318.170 ;
        RECT 268.340 33.310 268.480 1317.850 ;
        RECT 268.280 32.990 268.540 33.310 ;
        RECT 888.820 32.990 889.080 33.310 ;
        RECT 888.880 2.400 889.020 32.990 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 910.410 68.920 910.730 68.980 ;
        RECT 925.590 68.920 925.910 68.980 ;
        RECT 910.410 68.780 925.910 68.920 ;
        RECT 910.410 68.720 910.730 68.780 ;
        RECT 925.590 68.720 925.910 68.780 ;
        RECT 906.730 16.900 907.050 16.960 ;
        RECT 910.410 16.900 910.730 16.960 ;
        RECT 906.730 16.760 910.730 16.900 ;
        RECT 906.730 16.700 907.050 16.760 ;
        RECT 910.410 16.700 910.730 16.760 ;
      LAYER via ;
        RECT 910.440 68.720 910.700 68.980 ;
        RECT 925.620 68.720 925.880 68.980 ;
        RECT 906.760 16.700 907.020 16.960 ;
        RECT 910.440 16.700 910.700 16.960 ;
      LAYER met2 ;
        RECT 930.170 216.650 930.450 220.000 ;
        RECT 927.980 216.510 930.450 216.650 ;
        RECT 927.980 159.530 928.120 216.510 ;
        RECT 930.170 216.000 930.450 216.510 ;
        RECT 926.600 159.390 928.120 159.530 ;
        RECT 926.600 158.850 926.740 159.390 ;
        RECT 925.680 158.710 926.740 158.850 ;
        RECT 925.680 69.010 925.820 158.710 ;
        RECT 910.440 68.690 910.700 69.010 ;
        RECT 925.620 68.690 925.880 69.010 ;
        RECT 910.500 16.990 910.640 68.690 ;
        RECT 906.760 16.670 907.020 16.990 ;
        RECT 910.440 16.670 910.700 16.990 ;
        RECT 906.820 2.400 906.960 16.670 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 917.770 16.900 918.090 16.960 ;
        RECT 924.210 16.900 924.530 16.960 ;
        RECT 917.770 16.760 924.530 16.900 ;
        RECT 917.770 16.700 918.090 16.760 ;
        RECT 924.210 16.700 924.530 16.760 ;
      LAYER via ;
        RECT 917.800 16.700 918.060 16.960 ;
        RECT 924.240 16.700 924.500 16.960 ;
      LAYER met2 ;
        RECT 311.970 1028.995 312.250 1029.365 ;
        RECT 312.040 1007.605 312.180 1028.995 ;
        RECT 311.970 1007.235 312.250 1007.605 ;
        RECT 311.970 640.715 312.250 641.085 ;
        RECT 312.040 580.565 312.180 640.715 ;
        RECT 311.970 580.195 312.250 580.565 ;
        RECT 311.970 557.075 312.250 557.445 ;
        RECT 312.040 531.605 312.180 557.075 ;
        RECT 311.970 531.235 312.250 531.605 ;
        RECT 311.050 529.875 311.330 530.245 ;
        RECT 311.120 491.485 311.260 529.875 ;
        RECT 311.050 491.115 311.330 491.485 ;
        RECT 311.970 468.675 312.250 469.045 ;
        RECT 312.040 443.205 312.180 468.675 ;
        RECT 311.970 442.835 312.250 443.205 ;
        RECT 311.050 352.395 311.330 352.765 ;
        RECT 311.120 303.805 311.260 352.395 ;
        RECT 311.050 303.435 311.330 303.805 ;
        RECT 917.790 154.515 918.070 154.885 ;
        RECT 917.860 16.990 918.000 154.515 ;
        RECT 917.800 16.670 918.060 16.990 ;
        RECT 924.240 16.670 924.500 16.990 ;
        RECT 924.300 2.400 924.440 16.670 ;
        RECT 924.090 -4.800 924.650 2.400 ;
      LAYER via2 ;
        RECT 311.970 1029.040 312.250 1029.320 ;
        RECT 311.970 1007.280 312.250 1007.560 ;
        RECT 311.970 640.760 312.250 641.040 ;
        RECT 311.970 580.240 312.250 580.520 ;
        RECT 311.970 557.120 312.250 557.400 ;
        RECT 311.970 531.280 312.250 531.560 ;
        RECT 311.050 529.920 311.330 530.200 ;
        RECT 311.050 491.160 311.330 491.440 ;
        RECT 311.970 468.720 312.250 469.000 ;
        RECT 311.970 442.880 312.250 443.160 ;
        RECT 311.050 352.440 311.330 352.720 ;
        RECT 311.050 303.480 311.330 303.760 ;
        RECT 917.790 154.560 918.070 154.840 ;
      LAYER met3 ;
        RECT 310.000 1221.080 314.000 1221.680 ;
        RECT 313.110 1219.060 313.410 1221.080 ;
        RECT 313.070 1218.740 313.450 1219.060 ;
        RECT 311.945 1029.330 312.275 1029.345 ;
        RECT 313.070 1029.330 313.450 1029.340 ;
        RECT 311.945 1029.030 313.450 1029.330 ;
        RECT 311.945 1029.015 312.275 1029.030 ;
        RECT 313.070 1029.020 313.450 1029.030 ;
        RECT 311.945 1007.570 312.275 1007.585 ;
        RECT 313.070 1007.570 313.450 1007.580 ;
        RECT 311.945 1007.270 313.450 1007.570 ;
        RECT 311.945 1007.255 312.275 1007.270 ;
        RECT 313.070 1007.260 313.450 1007.270 ;
        RECT 313.070 919.170 313.450 919.180 ;
        RECT 312.190 918.870 313.450 919.170 ;
        RECT 312.190 918.500 312.490 918.870 ;
        RECT 313.070 918.860 313.450 918.870 ;
        RECT 312.150 918.180 312.530 918.500 ;
        RECT 310.310 772.970 310.690 772.980 ;
        RECT 312.150 772.970 312.530 772.980 ;
        RECT 310.310 772.670 312.530 772.970 ;
        RECT 310.310 772.660 310.690 772.670 ;
        RECT 312.150 772.660 312.530 772.670 ;
        RECT 310.310 718.260 310.690 718.580 ;
        RECT 310.350 717.890 310.650 718.260 ;
        RECT 313.070 717.890 313.450 717.900 ;
        RECT 310.350 717.590 313.450 717.890 ;
        RECT 313.070 717.580 313.450 717.590 ;
        RECT 311.230 641.050 311.610 641.060 ;
        RECT 311.945 641.050 312.275 641.065 ;
        RECT 311.230 640.750 312.275 641.050 ;
        RECT 311.230 640.740 311.610 640.750 ;
        RECT 311.945 640.735 312.275 640.750 ;
        RECT 311.945 580.530 312.275 580.545 ;
        RECT 311.945 580.215 312.490 580.530 ;
        RECT 312.190 579.860 312.490 580.215 ;
        RECT 312.150 579.540 312.530 579.860 ;
        RECT 311.945 557.410 312.275 557.425 ;
        RECT 313.070 557.410 313.450 557.420 ;
        RECT 311.945 557.110 313.450 557.410 ;
        RECT 311.945 557.095 312.275 557.110 ;
        RECT 313.070 557.100 313.450 557.110 ;
        RECT 311.945 531.570 312.275 531.585 ;
        RECT 313.070 531.570 313.450 531.580 ;
        RECT 311.945 531.270 313.450 531.570 ;
        RECT 311.945 531.255 312.275 531.270 ;
        RECT 313.070 531.260 313.450 531.270 ;
        RECT 311.025 530.210 311.355 530.225 ;
        RECT 313.070 530.210 313.450 530.220 ;
        RECT 311.025 529.910 313.450 530.210 ;
        RECT 311.025 529.895 311.355 529.910 ;
        RECT 313.070 529.900 313.450 529.910 ;
        RECT 311.025 491.450 311.355 491.465 ;
        RECT 313.070 491.450 313.450 491.460 ;
        RECT 311.025 491.150 313.450 491.450 ;
        RECT 311.025 491.135 311.355 491.150 ;
        RECT 313.070 491.140 313.450 491.150 ;
        RECT 311.945 469.010 312.275 469.025 ;
        RECT 313.070 469.010 313.450 469.020 ;
        RECT 311.945 468.710 313.450 469.010 ;
        RECT 311.945 468.695 312.275 468.710 ;
        RECT 313.070 468.700 313.450 468.710 ;
        RECT 311.945 443.170 312.275 443.185 ;
        RECT 313.070 443.170 313.450 443.180 ;
        RECT 311.945 442.870 313.450 443.170 ;
        RECT 311.945 442.855 312.275 442.870 ;
        RECT 313.070 442.860 313.450 442.870 ;
        RECT 311.025 352.730 311.355 352.745 ;
        RECT 313.070 352.730 313.450 352.740 ;
        RECT 311.025 352.430 313.450 352.730 ;
        RECT 311.025 352.415 311.355 352.430 ;
        RECT 313.070 352.420 313.450 352.430 ;
        RECT 311.025 303.770 311.355 303.785 ;
        RECT 313.070 303.770 313.450 303.780 ;
        RECT 311.025 303.470 313.450 303.770 ;
        RECT 311.025 303.455 311.355 303.470 ;
        RECT 313.070 303.460 313.450 303.470 ;
        RECT 310.310 262.290 310.690 262.300 ;
        RECT 313.070 262.290 313.450 262.300 ;
        RECT 310.310 261.990 313.450 262.290 ;
        RECT 310.310 261.980 310.690 261.990 ;
        RECT 313.070 261.980 313.450 261.990 ;
        RECT 310.310 218.770 310.690 218.780 ;
        RECT 313.990 218.770 314.370 218.780 ;
        RECT 310.310 218.470 314.370 218.770 ;
        RECT 310.310 218.460 310.690 218.470 ;
        RECT 313.990 218.460 314.370 218.470 ;
        RECT 313.070 154.850 313.450 154.860 ;
        RECT 917.765 154.850 918.095 154.865 ;
        RECT 313.070 154.550 918.095 154.850 ;
        RECT 313.070 154.540 313.450 154.550 ;
        RECT 917.765 154.535 918.095 154.550 ;
      LAYER via3 ;
        RECT 313.100 1218.740 313.420 1219.060 ;
        RECT 313.100 1029.020 313.420 1029.340 ;
        RECT 313.100 1007.260 313.420 1007.580 ;
        RECT 313.100 918.860 313.420 919.180 ;
        RECT 312.180 918.180 312.500 918.500 ;
        RECT 310.340 772.660 310.660 772.980 ;
        RECT 312.180 772.660 312.500 772.980 ;
        RECT 310.340 718.260 310.660 718.580 ;
        RECT 313.100 717.580 313.420 717.900 ;
        RECT 311.260 640.740 311.580 641.060 ;
        RECT 312.180 579.540 312.500 579.860 ;
        RECT 313.100 557.100 313.420 557.420 ;
        RECT 313.100 531.260 313.420 531.580 ;
        RECT 313.100 529.900 313.420 530.220 ;
        RECT 313.100 491.140 313.420 491.460 ;
        RECT 313.100 468.700 313.420 469.020 ;
        RECT 313.100 442.860 313.420 443.180 ;
        RECT 313.100 352.420 313.420 352.740 ;
        RECT 313.100 303.460 313.420 303.780 ;
        RECT 310.340 261.980 310.660 262.300 ;
        RECT 313.100 261.980 313.420 262.300 ;
        RECT 310.340 218.460 310.660 218.780 ;
        RECT 314.020 218.460 314.340 218.780 ;
        RECT 313.100 154.540 313.420 154.860 ;
      LAYER met4 ;
        RECT 313.095 1218.735 313.425 1219.065 ;
        RECT 313.110 1174.850 313.410 1218.735 ;
        RECT 312.190 1174.550 313.410 1174.850 ;
        RECT 312.190 1123.850 312.490 1174.550 ;
        RECT 312.190 1123.550 313.410 1123.850 ;
        RECT 313.110 1029.345 313.410 1123.550 ;
        RECT 313.095 1029.015 313.425 1029.345 ;
        RECT 313.095 1007.255 313.425 1007.585 ;
        RECT 313.110 919.185 313.410 1007.255 ;
        RECT 313.095 918.855 313.425 919.185 ;
        RECT 312.175 918.175 312.505 918.505 ;
        RECT 312.190 772.985 312.490 918.175 ;
        RECT 310.335 772.655 310.665 772.985 ;
        RECT 312.175 772.655 312.505 772.985 ;
        RECT 310.350 718.585 310.650 772.655 ;
        RECT 310.335 718.255 310.665 718.585 ;
        RECT 313.095 717.575 313.425 717.905 ;
        RECT 313.110 685.250 313.410 717.575 ;
        RECT 311.270 684.950 313.410 685.250 ;
        RECT 311.270 641.065 311.570 684.950 ;
        RECT 311.255 640.735 311.585 641.065 ;
        RECT 312.175 579.850 312.505 579.865 ;
        RECT 312.175 579.550 313.410 579.850 ;
        RECT 312.175 579.535 312.505 579.550 ;
        RECT 313.110 557.425 313.410 579.550 ;
        RECT 313.095 557.095 313.425 557.425 ;
        RECT 313.095 531.255 313.425 531.585 ;
        RECT 313.110 530.225 313.410 531.255 ;
        RECT 313.095 529.895 313.425 530.225 ;
        RECT 313.095 491.135 313.425 491.465 ;
        RECT 313.110 469.025 313.410 491.135 ;
        RECT 313.095 468.695 313.425 469.025 ;
        RECT 313.095 442.855 313.425 443.185 ;
        RECT 313.110 416.650 313.410 442.855 ;
        RECT 312.190 416.350 313.410 416.650 ;
        RECT 312.190 396.250 312.490 416.350 ;
        RECT 312.190 395.950 313.410 396.250 ;
        RECT 313.110 352.745 313.410 395.950 ;
        RECT 313.095 352.415 313.425 352.745 ;
        RECT 313.095 303.455 313.425 303.785 ;
        RECT 313.110 262.305 313.410 303.455 ;
        RECT 310.335 261.975 310.665 262.305 ;
        RECT 313.095 261.975 313.425 262.305 ;
        RECT 310.350 218.785 310.650 261.975 ;
        RECT 310.335 218.455 310.665 218.785 ;
        RECT 314.015 218.455 314.345 218.785 ;
        RECT 314.030 205.850 314.330 218.455 ;
        RECT 313.110 205.550 314.330 205.850 ;
        RECT 313.110 154.865 313.410 205.550 ;
        RECT 313.095 154.535 313.425 154.865 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 306.430 218.520 306.750 218.580 ;
        RECT 938.470 218.520 938.790 218.580 ;
        RECT 306.430 218.380 938.790 218.520 ;
        RECT 306.430 218.320 306.750 218.380 ;
        RECT 938.470 218.320 938.790 218.380 ;
        RECT 938.470 2.960 938.790 3.020 ;
        RECT 942.150 2.960 942.470 3.020 ;
        RECT 938.470 2.820 942.470 2.960 ;
        RECT 938.470 2.760 938.790 2.820 ;
        RECT 942.150 2.760 942.470 2.820 ;
      LAYER via ;
        RECT 306.460 218.320 306.720 218.580 ;
        RECT 938.500 218.320 938.760 218.580 ;
        RECT 938.500 2.760 938.760 3.020 ;
        RECT 942.180 2.760 942.440 3.020 ;
      LAYER met2 ;
        RECT 306.450 957.595 306.730 957.965 ;
        RECT 306.520 218.610 306.660 957.595 ;
        RECT 306.460 218.290 306.720 218.610 ;
        RECT 938.500 218.290 938.760 218.610 ;
        RECT 938.560 3.050 938.700 218.290 ;
        RECT 938.500 2.730 938.760 3.050 ;
        RECT 942.180 2.730 942.440 3.050 ;
        RECT 942.240 2.400 942.380 2.730 ;
        RECT 942.030 -4.800 942.590 2.400 ;
      LAYER via2 ;
        RECT 306.450 957.640 306.730 957.920 ;
      LAYER met3 ;
        RECT 306.425 957.930 306.755 957.945 ;
        RECT 306.425 957.840 310.500 957.930 ;
        RECT 306.425 957.630 314.000 957.840 ;
        RECT 306.425 957.615 306.755 957.630 ;
        RECT 310.000 957.240 314.000 957.630 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.950 1342.220 864.270 1342.280 ;
        RECT 1409.050 1342.220 1409.370 1342.280 ;
        RECT 863.950 1342.080 1409.370 1342.220 ;
        RECT 863.950 1342.020 864.270 1342.080 ;
        RECT 1409.050 1342.020 1409.370 1342.080 ;
        RECT 960.090 33.900 960.410 33.960 ;
        RECT 1409.050 33.900 1409.370 33.960 ;
        RECT 960.090 33.760 1409.370 33.900 ;
        RECT 960.090 33.700 960.410 33.760 ;
        RECT 1409.050 33.700 1409.370 33.760 ;
      LAYER via ;
        RECT 863.980 1342.020 864.240 1342.280 ;
        RECT 1409.080 1342.020 1409.340 1342.280 ;
        RECT 960.120 33.700 960.380 33.960 ;
        RECT 1409.080 33.700 1409.340 33.960 ;
      LAYER met2 ;
        RECT 863.980 1341.990 864.240 1342.310 ;
        RECT 1409.080 1341.990 1409.340 1342.310 ;
        RECT 864.040 1325.025 864.180 1341.990 ;
        RECT 863.930 1321.025 864.210 1325.025 ;
        RECT 1409.140 33.990 1409.280 1341.990 ;
        RECT 960.120 33.670 960.380 33.990 ;
        RECT 1409.080 33.670 1409.340 33.990 ;
        RECT 960.180 2.400 960.320 33.670 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 268.710 1332.020 269.030 1332.080 ;
        RECT 329.430 1332.020 329.750 1332.080 ;
        RECT 268.710 1331.880 329.750 1332.020 ;
        RECT 268.710 1331.820 269.030 1331.880 ;
        RECT 329.430 1331.820 329.750 1331.880 ;
        RECT 268.710 32.200 269.030 32.260 ;
        RECT 978.030 32.200 978.350 32.260 ;
        RECT 268.710 32.060 978.350 32.200 ;
        RECT 268.710 32.000 269.030 32.060 ;
        RECT 978.030 32.000 978.350 32.060 ;
      LAYER via ;
        RECT 268.740 1331.820 269.000 1332.080 ;
        RECT 329.460 1331.820 329.720 1332.080 ;
        RECT 268.740 32.000 269.000 32.260 ;
        RECT 978.060 32.000 978.320 32.260 ;
      LAYER met2 ;
        RECT 268.740 1331.790 269.000 1332.110 ;
        RECT 329.460 1331.790 329.720 1332.110 ;
        RECT 268.800 32.290 268.940 1331.790 ;
        RECT 329.520 1325.025 329.660 1331.790 ;
        RECT 329.410 1321.025 329.690 1325.025 ;
        RECT 268.740 31.970 269.000 32.290 ;
        RECT 978.060 31.970 978.320 32.290 ;
        RECT 978.120 2.400 978.260 31.970 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.950 59.740 657.270 59.800 ;
        RECT 1409.510 59.740 1409.830 59.800 ;
        RECT 656.950 59.600 1409.830 59.740 ;
        RECT 656.950 59.540 657.270 59.600 ;
        RECT 1409.510 59.540 1409.830 59.600 ;
      LAYER via ;
        RECT 656.980 59.540 657.240 59.800 ;
        RECT 1409.540 59.540 1409.800 59.800 ;
      LAYER met2 ;
        RECT 1409.530 314.315 1409.810 314.685 ;
        RECT 1409.600 59.830 1409.740 314.315 ;
        RECT 656.980 59.510 657.240 59.830 ;
        RECT 1409.540 59.510 1409.800 59.830 ;
        RECT 657.040 2.400 657.180 59.510 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 1409.530 314.360 1409.810 314.640 ;
      LAYER met3 ;
        RECT 1409.505 314.650 1409.835 314.665 ;
        RECT 1408.060 314.560 1409.835 314.650 ;
        RECT 1404.305 314.350 1409.835 314.560 ;
        RECT 1404.305 313.960 1408.305 314.350 ;
        RECT 1409.505 314.335 1409.835 314.350 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1185.030 1334.740 1185.350 1334.800 ;
        RECT 1408.590 1334.740 1408.910 1334.800 ;
        RECT 1185.030 1334.600 1408.910 1334.740 ;
        RECT 1185.030 1334.540 1185.350 1334.600 ;
        RECT 1408.590 1334.540 1408.910 1334.600 ;
        RECT 995.970 19.620 996.290 19.680 ;
        RECT 1408.590 19.620 1408.910 19.680 ;
        RECT 995.970 19.480 1408.910 19.620 ;
        RECT 995.970 19.420 996.290 19.480 ;
        RECT 1408.590 19.420 1408.910 19.480 ;
      LAYER via ;
        RECT 1185.060 1334.540 1185.320 1334.800 ;
        RECT 1408.620 1334.540 1408.880 1334.800 ;
        RECT 996.000 19.420 996.260 19.680 ;
        RECT 1408.620 19.420 1408.880 19.680 ;
      LAYER met2 ;
        RECT 1185.060 1334.510 1185.320 1334.830 ;
        RECT 1408.620 1334.510 1408.880 1334.830 ;
        RECT 1185.120 1325.025 1185.260 1334.510 ;
        RECT 1185.010 1321.025 1185.290 1325.025 ;
        RECT 1408.680 19.710 1408.820 1334.510 ;
        RECT 996.000 19.390 996.260 19.710 ;
        RECT 1408.620 19.390 1408.880 19.710 ;
        RECT 996.060 2.400 996.200 19.390 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1405.370 190.300 1405.690 190.360 ;
        RECT 1393.040 190.160 1405.690 190.300 ;
        RECT 1013.910 189.960 1014.230 190.020 ;
        RECT 1393.040 189.960 1393.180 190.160 ;
        RECT 1405.370 190.100 1405.690 190.160 ;
        RECT 1013.910 189.820 1393.180 189.960 ;
        RECT 1013.910 189.760 1014.230 189.820 ;
      LAYER via ;
        RECT 1013.940 189.760 1014.200 190.020 ;
        RECT 1405.400 190.100 1405.660 190.360 ;
      LAYER met2 ;
        RECT 1405.390 297.995 1405.670 298.365 ;
        RECT 1405.460 190.390 1405.600 297.995 ;
        RECT 1405.400 190.070 1405.660 190.390 ;
        RECT 1013.940 189.730 1014.200 190.050 ;
        RECT 1014.000 17.410 1014.140 189.730 ;
        RECT 1013.540 17.270 1014.140 17.410 ;
        RECT 1013.540 2.400 1013.680 17.270 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
      LAYER via2 ;
        RECT 1405.390 298.040 1405.670 298.320 ;
      LAYER met3 ;
        RECT 1404.305 300.360 1408.305 300.960 ;
        RECT 1405.150 298.345 1405.450 300.360 ;
        RECT 1405.150 298.030 1405.695 298.345 ;
        RECT 1405.365 298.015 1405.695 298.030 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 301.830 214.780 302.150 214.840 ;
        RECT 320.690 214.780 321.010 214.840 ;
        RECT 301.830 214.640 321.010 214.780 ;
        RECT 301.830 214.580 302.150 214.640 ;
        RECT 320.690 214.580 321.010 214.640 ;
        RECT 320.690 17.920 321.010 17.980 ;
        RECT 1031.390 17.920 1031.710 17.980 ;
        RECT 320.690 17.780 1031.710 17.920 ;
        RECT 320.690 17.720 321.010 17.780 ;
        RECT 1031.390 17.720 1031.710 17.780 ;
      LAYER via ;
        RECT 301.860 214.580 302.120 214.840 ;
        RECT 320.720 214.580 320.980 214.840 ;
        RECT 320.720 17.720 320.980 17.980 ;
        RECT 1031.420 17.720 1031.680 17.980 ;
      LAYER met2 ;
        RECT 301.850 965.755 302.130 966.125 ;
        RECT 301.920 214.870 302.060 965.755 ;
        RECT 301.860 214.550 302.120 214.870 ;
        RECT 320.720 214.550 320.980 214.870 ;
        RECT 320.780 18.010 320.920 214.550 ;
        RECT 320.720 17.690 320.980 18.010 ;
        RECT 1031.420 17.690 1031.680 18.010 ;
        RECT 1031.480 2.400 1031.620 17.690 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
      LAYER via2 ;
        RECT 301.850 965.800 302.130 966.080 ;
      LAYER met3 ;
        RECT 301.825 966.090 302.155 966.105 ;
        RECT 301.825 966.000 310.500 966.090 ;
        RECT 301.825 965.790 314.000 966.000 ;
        RECT 301.825 965.775 302.155 965.790 ;
        RECT 310.000 965.400 314.000 965.790 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.450 1321.650 1007.730 1325.025 ;
        RECT 1008.410 1321.650 1008.690 1321.765 ;
        RECT 1007.450 1321.510 1008.690 1321.650 ;
        RECT 1007.450 1321.025 1007.730 1321.510 ;
        RECT 1008.410 1321.395 1008.690 1321.510 ;
        RECT 1049.350 30.075 1049.630 30.445 ;
        RECT 1049.420 2.400 1049.560 30.075 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
      LAYER via2 ;
        RECT 1008.410 1321.440 1008.690 1321.720 ;
        RECT 1049.350 30.120 1049.630 30.400 ;
      LAYER met3 ;
        RECT 1008.385 1321.740 1008.715 1321.745 ;
        RECT 1008.385 1321.730 1008.970 1321.740 ;
        RECT 1008.385 1321.430 1009.170 1321.730 ;
        RECT 1008.385 1321.420 1008.970 1321.430 ;
        RECT 1008.385 1321.415 1008.715 1321.420 ;
        RECT 1049.325 30.410 1049.655 30.425 ;
        RECT 1421.670 30.410 1422.050 30.420 ;
        RECT 1049.325 30.110 1422.050 30.410 ;
        RECT 1049.325 30.095 1049.655 30.110 ;
        RECT 1421.670 30.100 1422.050 30.110 ;
      LAYER via3 ;
        RECT 1008.620 1321.420 1008.940 1321.740 ;
        RECT 1421.700 30.100 1422.020 30.420 ;
      LAYER met4 ;
        RECT 1008.615 1321.415 1008.945 1321.745 ;
        RECT 1008.630 1314.690 1008.930 1321.415 ;
        RECT 1008.190 1313.510 1009.370 1314.690 ;
        RECT 1421.270 1313.510 1422.450 1314.690 ;
        RECT 1421.710 30.425 1422.010 1313.510 ;
        RECT 1421.695 30.095 1422.025 30.425 ;
      LAYER met5 ;
        RECT 1007.980 1313.300 1422.660 1314.900 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 274.690 1069.880 275.010 1069.940 ;
        RECT 296.770 1069.880 297.090 1069.940 ;
        RECT 274.690 1069.740 297.090 1069.880 ;
        RECT 274.690 1069.680 275.010 1069.740 ;
        RECT 296.770 1069.680 297.090 1069.740 ;
        RECT 274.690 31.180 275.010 31.240 ;
        RECT 1067.270 31.180 1067.590 31.240 ;
        RECT 274.690 31.040 1067.590 31.180 ;
        RECT 274.690 30.980 275.010 31.040 ;
        RECT 1067.270 30.980 1067.590 31.040 ;
      LAYER via ;
        RECT 274.720 1069.680 274.980 1069.940 ;
        RECT 296.800 1069.680 297.060 1069.940 ;
        RECT 274.720 30.980 274.980 31.240 ;
        RECT 1067.300 30.980 1067.560 31.240 ;
      LAYER met2 ;
        RECT 296.790 1074.555 297.070 1074.925 ;
        RECT 296.860 1069.970 297.000 1074.555 ;
        RECT 274.720 1069.650 274.980 1069.970 ;
        RECT 296.800 1069.650 297.060 1069.970 ;
        RECT 274.780 31.270 274.920 1069.650 ;
        RECT 274.720 30.950 274.980 31.270 ;
        RECT 1067.300 30.950 1067.560 31.270 ;
        RECT 1067.360 2.400 1067.500 30.950 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
      LAYER via2 ;
        RECT 296.790 1074.600 297.070 1074.880 ;
      LAYER met3 ;
        RECT 296.765 1074.890 297.095 1074.905 ;
        RECT 296.765 1074.800 310.500 1074.890 ;
        RECT 296.765 1074.590 314.000 1074.800 ;
        RECT 296.765 1074.575 297.095 1074.590 ;
        RECT 310.000 1074.200 314.000 1074.590 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1210.790 135.220 1211.110 135.280 ;
        RECT 1419.630 135.220 1419.950 135.280 ;
        RECT 1210.790 135.080 1419.950 135.220 ;
        RECT 1210.790 135.020 1211.110 135.080 ;
        RECT 1419.630 135.020 1419.950 135.080 ;
        RECT 1085.210 19.280 1085.530 19.340 ;
        RECT 1210.790 19.280 1211.110 19.340 ;
        RECT 1085.210 19.140 1211.110 19.280 ;
        RECT 1085.210 19.080 1085.530 19.140 ;
        RECT 1210.790 19.080 1211.110 19.140 ;
      LAYER via ;
        RECT 1210.820 135.020 1211.080 135.280 ;
        RECT 1419.660 135.020 1419.920 135.280 ;
        RECT 1085.240 19.080 1085.500 19.340 ;
        RECT 1210.820 19.080 1211.080 19.340 ;
      LAYER met2 ;
        RECT 1419.650 922.235 1419.930 922.605 ;
        RECT 1419.720 135.310 1419.860 922.235 ;
        RECT 1210.820 134.990 1211.080 135.310 ;
        RECT 1419.660 134.990 1419.920 135.310 ;
        RECT 1210.880 19.370 1211.020 134.990 ;
        RECT 1085.240 19.050 1085.500 19.370 ;
        RECT 1210.820 19.050 1211.080 19.370 ;
        RECT 1085.300 2.400 1085.440 19.050 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
      LAYER via2 ;
        RECT 1419.650 922.280 1419.930 922.560 ;
      LAYER met3 ;
        RECT 1419.625 922.570 1419.955 922.585 ;
        RECT 1408.060 922.480 1419.955 922.570 ;
        RECT 1404.305 922.270 1419.955 922.480 ;
        RECT 1404.305 921.880 1408.305 922.270 ;
        RECT 1419.625 922.255 1419.955 922.270 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1103.610 122.300 1103.930 122.360 ;
        RECT 1415.030 122.300 1415.350 122.360 ;
        RECT 1103.610 122.160 1415.350 122.300 ;
        RECT 1103.610 122.100 1103.930 122.160 ;
        RECT 1415.030 122.100 1415.350 122.160 ;
      LAYER via ;
        RECT 1103.640 122.100 1103.900 122.360 ;
        RECT 1415.060 122.100 1415.320 122.360 ;
      LAYER met2 ;
        RECT 1415.050 965.755 1415.330 966.125 ;
        RECT 1415.120 122.390 1415.260 965.755 ;
        RECT 1103.640 122.070 1103.900 122.390 ;
        RECT 1415.060 122.070 1415.320 122.390 ;
        RECT 1103.700 17.410 1103.840 122.070 ;
        RECT 1102.780 17.270 1103.840 17.410 ;
        RECT 1102.780 2.400 1102.920 17.270 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
      LAYER via2 ;
        RECT 1415.050 965.800 1415.330 966.080 ;
      LAYER met3 ;
        RECT 1415.025 966.090 1415.355 966.105 ;
        RECT 1408.060 966.000 1415.355 966.090 ;
        RECT 1404.305 965.790 1415.355 966.000 ;
        RECT 1404.305 965.400 1408.305 965.790 ;
        RECT 1415.025 965.775 1415.355 965.790 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 310.110 218.180 310.430 218.240 ;
        RECT 1119.250 218.180 1119.570 218.240 ;
        RECT 310.110 218.040 1119.570 218.180 ;
        RECT 310.110 217.980 310.430 218.040 ;
        RECT 1119.250 217.980 1119.570 218.040 ;
      LAYER via ;
        RECT 310.140 217.980 310.400 218.240 ;
        RECT 1119.280 217.980 1119.540 218.240 ;
      LAYER met2 ;
        RECT 310.130 231.355 310.410 231.725 ;
        RECT 310.200 218.270 310.340 231.355 ;
        RECT 310.140 217.950 310.400 218.270 ;
        RECT 1119.280 217.950 1119.540 218.270 ;
        RECT 1119.340 17.410 1119.480 217.950 ;
        RECT 1119.340 17.270 1120.860 17.410 ;
        RECT 1120.720 2.400 1120.860 17.270 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
      LAYER via2 ;
        RECT 310.130 231.400 310.410 231.680 ;
      LAYER met3 ;
        RECT 310.000 233.720 314.000 234.320 ;
        RECT 310.350 231.705 310.650 233.720 ;
        RECT 310.105 231.390 310.650 231.705 ;
        RECT 310.105 231.375 310.435 231.390 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 299.990 217.840 300.310 217.900 ;
        RECT 1138.570 217.840 1138.890 217.900 ;
        RECT 299.990 217.700 1138.890 217.840 ;
        RECT 299.990 217.640 300.310 217.700 ;
        RECT 1138.570 217.640 1138.890 217.700 ;
      LAYER via ;
        RECT 300.020 217.640 300.280 217.900 ;
        RECT 1138.600 217.640 1138.860 217.900 ;
      LAYER met2 ;
        RECT 300.010 402.715 300.290 403.085 ;
        RECT 300.080 217.930 300.220 402.715 ;
        RECT 300.020 217.610 300.280 217.930 ;
        RECT 1138.600 217.610 1138.860 217.930 ;
        RECT 1138.660 2.400 1138.800 217.610 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
      LAYER via2 ;
        RECT 300.010 402.760 300.290 403.040 ;
      LAYER met3 ;
        RECT 299.985 403.050 300.315 403.065 ;
        RECT 299.985 402.960 310.500 403.050 ;
        RECT 299.985 402.750 314.000 402.960 ;
        RECT 299.985 402.735 300.315 402.750 ;
        RECT 310.000 402.360 314.000 402.750 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1158.810 80.820 1159.130 80.880 ;
        RECT 1417.790 80.820 1418.110 80.880 ;
        RECT 1158.810 80.680 1418.110 80.820 ;
        RECT 1158.810 80.620 1159.130 80.680 ;
        RECT 1417.790 80.620 1418.110 80.680 ;
        RECT 1156.510 16.900 1156.830 16.960 ;
        RECT 1158.810 16.900 1159.130 16.960 ;
        RECT 1156.510 16.760 1159.130 16.900 ;
        RECT 1156.510 16.700 1156.830 16.760 ;
        RECT 1158.810 16.700 1159.130 16.760 ;
      LAYER via ;
        RECT 1158.840 80.620 1159.100 80.880 ;
        RECT 1417.820 80.620 1418.080 80.880 ;
        RECT 1156.540 16.700 1156.800 16.960 ;
        RECT 1158.840 16.700 1159.100 16.960 ;
      LAYER met2 ;
        RECT 1417.810 584.955 1418.090 585.325 ;
        RECT 1417.880 80.910 1418.020 584.955 ;
        RECT 1158.840 80.590 1159.100 80.910 ;
        RECT 1417.820 80.590 1418.080 80.910 ;
        RECT 1158.900 16.990 1159.040 80.590 ;
        RECT 1156.540 16.670 1156.800 16.990 ;
        RECT 1158.840 16.670 1159.100 16.990 ;
        RECT 1156.600 2.400 1156.740 16.670 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
      LAYER via2 ;
        RECT 1417.810 585.000 1418.090 585.280 ;
      LAYER met3 ;
        RECT 1417.785 585.290 1418.115 585.305 ;
        RECT 1408.060 585.200 1418.115 585.290 ;
        RECT 1404.305 584.990 1418.115 585.200 ;
        RECT 1404.305 584.600 1408.305 584.990 ;
        RECT 1417.785 584.975 1418.115 584.990 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 675.425 193.205 675.595 210.715 ;
        RECT 675.425 144.925 675.595 192.695 ;
        RECT 675.885 48.365 676.055 96.135 ;
      LAYER mcon ;
        RECT 675.425 210.545 675.595 210.715 ;
        RECT 675.425 192.525 675.595 192.695 ;
        RECT 675.885 95.965 676.055 96.135 ;
      LAYER met1 ;
        RECT 1303.710 1345.620 1304.030 1345.680 ;
        RECT 1430.210 1345.620 1430.530 1345.680 ;
        RECT 1303.710 1345.480 1430.530 1345.620 ;
        RECT 1303.710 1345.420 1304.030 1345.480 ;
        RECT 1430.210 1345.420 1430.530 1345.480 ;
        RECT 675.365 210.700 675.655 210.745 ;
        RECT 1430.210 210.700 1430.530 210.760 ;
        RECT 675.365 210.560 1430.530 210.700 ;
        RECT 675.365 210.515 675.655 210.560 ;
        RECT 1430.210 210.500 1430.530 210.560 ;
        RECT 675.365 193.360 675.655 193.405 ;
        RECT 675.810 193.360 676.130 193.420 ;
        RECT 675.365 193.220 676.130 193.360 ;
        RECT 675.365 193.175 675.655 193.220 ;
        RECT 675.810 193.160 676.130 193.220 ;
        RECT 675.365 192.680 675.655 192.725 ;
        RECT 675.810 192.680 676.130 192.740 ;
        RECT 675.365 192.540 676.130 192.680 ;
        RECT 675.365 192.495 675.655 192.540 ;
        RECT 675.810 192.480 676.130 192.540 ;
        RECT 675.365 145.080 675.655 145.125 ;
        RECT 675.810 145.080 676.130 145.140 ;
        RECT 675.365 144.940 676.130 145.080 ;
        RECT 675.365 144.895 675.655 144.940 ;
        RECT 675.810 144.880 676.130 144.940 ;
        RECT 675.810 97.960 676.130 98.220 ;
        RECT 675.900 96.860 676.040 97.960 ;
        RECT 675.810 96.600 676.130 96.860 ;
        RECT 675.810 96.120 676.130 96.180 ;
        RECT 675.615 95.980 676.130 96.120 ;
        RECT 675.810 95.920 676.130 95.980 ;
        RECT 674.430 48.520 674.750 48.580 ;
        RECT 675.825 48.520 676.115 48.565 ;
        RECT 674.430 48.380 676.115 48.520 ;
        RECT 674.430 48.320 674.750 48.380 ;
        RECT 675.825 48.335 676.115 48.380 ;
      LAYER via ;
        RECT 1303.740 1345.420 1304.000 1345.680 ;
        RECT 1430.240 1345.420 1430.500 1345.680 ;
        RECT 1430.240 210.500 1430.500 210.760 ;
        RECT 675.840 193.160 676.100 193.420 ;
        RECT 675.840 192.480 676.100 192.740 ;
        RECT 675.840 144.880 676.100 145.140 ;
        RECT 675.840 97.960 676.100 98.220 ;
        RECT 675.840 96.600 676.100 96.860 ;
        RECT 675.840 95.920 676.100 96.180 ;
        RECT 674.460 48.320 674.720 48.580 ;
      LAYER met2 ;
        RECT 1303.740 1345.390 1304.000 1345.710 ;
        RECT 1430.240 1345.390 1430.500 1345.710 ;
        RECT 1303.800 1325.025 1303.940 1345.390 ;
        RECT 1303.690 1321.025 1303.970 1325.025 ;
        RECT 1430.300 210.790 1430.440 1345.390 ;
        RECT 1430.240 210.470 1430.500 210.790 ;
        RECT 675.840 193.130 676.100 193.450 ;
        RECT 675.900 192.770 676.040 193.130 ;
        RECT 675.840 192.450 676.100 192.770 ;
        RECT 675.840 144.850 676.100 145.170 ;
        RECT 675.900 98.250 676.040 144.850 ;
        RECT 675.840 97.930 676.100 98.250 ;
        RECT 675.840 96.570 676.100 96.890 ;
        RECT 675.900 96.210 676.040 96.570 ;
        RECT 675.840 95.890 676.100 96.210 ;
        RECT 674.460 48.290 674.720 48.610 ;
        RECT 674.520 2.400 674.660 48.290 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 620.610 142.700 620.930 142.760 ;
        RECT 1173.070 142.700 1173.390 142.760 ;
        RECT 620.610 142.560 1173.390 142.700 ;
        RECT 620.610 142.500 620.930 142.560 ;
        RECT 1173.070 142.500 1173.390 142.560 ;
        RECT 1172.610 48.520 1172.930 48.580 ;
        RECT 1173.990 48.520 1174.310 48.580 ;
        RECT 1172.610 48.380 1174.310 48.520 ;
        RECT 1172.610 48.320 1172.930 48.380 ;
        RECT 1173.990 48.320 1174.310 48.380 ;
      LAYER via ;
        RECT 620.640 142.500 620.900 142.760 ;
        RECT 1173.100 142.500 1173.360 142.760 ;
        RECT 1172.640 48.320 1172.900 48.580 ;
        RECT 1174.020 48.320 1174.280 48.580 ;
      LAYER met2 ;
        RECT 619.210 216.650 619.490 220.000 ;
        RECT 619.210 216.510 620.840 216.650 ;
        RECT 619.210 216.000 619.490 216.510 ;
        RECT 620.700 142.790 620.840 216.510 ;
        RECT 620.640 142.470 620.900 142.790 ;
        RECT 1173.100 142.470 1173.360 142.790 ;
        RECT 1173.160 72.490 1173.300 142.470 ;
        RECT 1172.700 72.350 1173.300 72.490 ;
        RECT 1172.700 48.610 1172.840 72.350 ;
        RECT 1172.640 48.290 1172.900 48.610 ;
        RECT 1174.020 48.290 1174.280 48.610 ;
        RECT 1174.080 2.400 1174.220 48.290 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 644.070 204.920 644.390 204.980 ;
        RECT 648.210 204.920 648.530 204.980 ;
        RECT 644.070 204.780 648.530 204.920 ;
        RECT 644.070 204.720 644.390 204.780 ;
        RECT 648.210 204.720 648.530 204.780 ;
        RECT 648.210 94.420 648.530 94.480 ;
        RECT 1187.790 94.420 1188.110 94.480 ;
        RECT 648.210 94.280 1188.110 94.420 ;
        RECT 648.210 94.220 648.530 94.280 ;
        RECT 1187.790 94.220 1188.110 94.280 ;
        RECT 1187.790 2.960 1188.110 3.020 ;
        RECT 1191.930 2.960 1192.250 3.020 ;
        RECT 1187.790 2.820 1192.250 2.960 ;
        RECT 1187.790 2.760 1188.110 2.820 ;
        RECT 1191.930 2.760 1192.250 2.820 ;
      LAYER via ;
        RECT 644.100 204.720 644.360 204.980 ;
        RECT 648.240 204.720 648.500 204.980 ;
        RECT 648.240 94.220 648.500 94.480 ;
        RECT 1187.820 94.220 1188.080 94.480 ;
        RECT 1187.820 2.760 1188.080 3.020 ;
        RECT 1191.960 2.760 1192.220 3.020 ;
      LAYER met2 ;
        RECT 644.050 216.000 644.330 220.000 ;
        RECT 644.160 205.010 644.300 216.000 ;
        RECT 644.100 204.690 644.360 205.010 ;
        RECT 648.240 204.690 648.500 205.010 ;
        RECT 648.300 94.510 648.440 204.690 ;
        RECT 648.240 94.190 648.500 94.510 ;
        RECT 1187.820 94.190 1188.080 94.510 ;
        RECT 1187.880 3.050 1188.020 94.190 ;
        RECT 1187.820 2.730 1188.080 3.050 ;
        RECT 1191.960 2.730 1192.220 3.050 ;
        RECT 1192.020 2.400 1192.160 2.730 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1209.870 25.740 1210.190 25.800 ;
        RECT 1418.250 25.740 1418.570 25.800 ;
        RECT 1209.870 25.600 1418.570 25.740 ;
        RECT 1209.870 25.540 1210.190 25.600 ;
        RECT 1418.250 25.540 1418.570 25.600 ;
      LAYER via ;
        RECT 1209.900 25.540 1210.160 25.800 ;
        RECT 1418.280 25.540 1418.540 25.800 ;
      LAYER met2 ;
        RECT 1418.270 402.715 1418.550 403.085 ;
        RECT 1418.340 25.830 1418.480 402.715 ;
        RECT 1209.900 25.510 1210.160 25.830 ;
        RECT 1418.280 25.510 1418.540 25.830 ;
        RECT 1209.960 2.400 1210.100 25.510 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
      LAYER via2 ;
        RECT 1418.270 402.760 1418.550 403.040 ;
      LAYER met3 ;
        RECT 1418.245 403.050 1418.575 403.065 ;
        RECT 1408.060 402.960 1418.575 403.050 ;
        RECT 1404.305 402.750 1418.575 402.960 ;
        RECT 1404.305 402.360 1408.305 402.750 ;
        RECT 1418.245 402.735 1418.575 402.750 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1415.950 190.980 1416.270 191.040 ;
        RECT 1392.120 190.840 1416.270 190.980 ;
        RECT 1227.810 190.640 1228.130 190.700 ;
        RECT 1392.120 190.640 1392.260 190.840 ;
        RECT 1415.950 190.780 1416.270 190.840 ;
        RECT 1227.810 190.500 1392.260 190.640 ;
        RECT 1227.810 190.440 1228.130 190.500 ;
      LAYER via ;
        RECT 1227.840 190.440 1228.100 190.700 ;
        RECT 1415.980 190.780 1416.240 191.040 ;
      LAYER met2 ;
        RECT 1416.430 263.995 1416.710 264.365 ;
        RECT 1416.500 245.890 1416.640 263.995 ;
        RECT 1416.040 245.750 1416.640 245.890 ;
        RECT 1416.040 191.070 1416.180 245.750 ;
        RECT 1415.980 190.750 1416.240 191.070 ;
        RECT 1227.840 190.410 1228.100 190.730 ;
        RECT 1227.900 2.400 1228.040 190.410 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
      LAYER via2 ;
        RECT 1416.430 264.040 1416.710 264.320 ;
      LAYER met3 ;
        RECT 1416.405 264.330 1416.735 264.345 ;
        RECT 1408.060 264.240 1416.735 264.330 ;
        RECT 1404.305 264.030 1416.735 264.240 ;
        RECT 1404.305 263.640 1408.305 264.030 ;
        RECT 1416.405 264.015 1416.735 264.030 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 344.610 114.820 344.930 114.880 ;
        RECT 1242.070 114.820 1242.390 114.880 ;
        RECT 344.610 114.680 1242.390 114.820 ;
        RECT 344.610 114.620 344.930 114.680 ;
        RECT 1242.070 114.620 1242.390 114.680 ;
      LAYER via ;
        RECT 344.640 114.620 344.900 114.880 ;
        RECT 1242.100 114.620 1242.360 114.880 ;
      LAYER met2 ;
        RECT 342.290 216.650 342.570 220.000 ;
        RECT 342.290 216.510 344.840 216.650 ;
        RECT 342.290 216.000 342.570 216.510 ;
        RECT 344.700 114.910 344.840 216.510 ;
        RECT 344.640 114.590 344.900 114.910 ;
        RECT 1242.100 114.590 1242.360 114.910 ;
        RECT 1242.160 17.410 1242.300 114.590 ;
        RECT 1242.160 17.270 1245.980 17.410 ;
        RECT 1245.840 2.400 1245.980 17.270 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 696.050 107.680 696.370 107.740 ;
        RECT 1263.230 107.680 1263.550 107.740 ;
        RECT 696.050 107.540 1263.550 107.680 ;
        RECT 696.050 107.480 696.370 107.540 ;
        RECT 1263.230 107.480 1263.550 107.540 ;
      LAYER via ;
        RECT 696.080 107.480 696.340 107.740 ;
        RECT 1263.260 107.480 1263.520 107.740 ;
      LAYER met2 ;
        RECT 692.810 216.650 693.090 220.000 ;
        RECT 692.810 216.510 696.280 216.650 ;
        RECT 692.810 216.000 693.090 216.510 ;
        RECT 696.140 107.770 696.280 216.510 ;
        RECT 696.080 107.450 696.340 107.770 ;
        RECT 1263.260 107.450 1263.520 107.770 ;
        RECT 1263.320 2.400 1263.460 107.450 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1282.550 66.200 1282.870 66.260 ;
        RECT 1416.870 66.200 1417.190 66.260 ;
        RECT 1282.550 66.060 1417.190 66.200 ;
        RECT 1282.550 66.000 1282.870 66.060 ;
        RECT 1416.870 66.000 1417.190 66.060 ;
      LAYER via ;
        RECT 1282.580 66.000 1282.840 66.260 ;
        RECT 1416.900 66.000 1417.160 66.260 ;
      LAYER met2 ;
        RECT 1416.890 629.835 1417.170 630.205 ;
        RECT 1416.960 66.290 1417.100 629.835 ;
        RECT 1282.580 65.970 1282.840 66.290 ;
        RECT 1416.900 65.970 1417.160 66.290 ;
        RECT 1282.640 17.410 1282.780 65.970 ;
        RECT 1281.260 17.270 1282.780 17.410 ;
        RECT 1281.260 2.400 1281.400 17.270 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
      LAYER via2 ;
        RECT 1416.890 629.880 1417.170 630.160 ;
      LAYER met3 ;
        RECT 1416.865 630.170 1417.195 630.185 ;
        RECT 1408.060 630.080 1417.195 630.170 ;
        RECT 1404.305 629.870 1417.195 630.080 ;
        RECT 1404.305 629.480 1408.305 629.870 ;
        RECT 1416.865 629.855 1417.195 629.870 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1261.005 1315.205 1261.175 1322.855 ;
      LAYER mcon ;
        RECT 1261.005 1322.685 1261.175 1322.855 ;
      LAYER met1 ;
        RECT 1260.930 1322.840 1261.250 1322.900 ;
        RECT 1260.735 1322.700 1261.250 1322.840 ;
        RECT 1260.930 1322.640 1261.250 1322.700 ;
        RECT 1260.945 1315.360 1261.235 1315.405 ;
        RECT 1429.290 1315.360 1429.610 1315.420 ;
        RECT 1260.945 1315.220 1429.610 1315.360 ;
        RECT 1260.945 1315.175 1261.235 1315.220 ;
        RECT 1429.290 1315.160 1429.610 1315.220 ;
        RECT 1299.110 16.560 1299.430 16.620 ;
        RECT 1429.290 16.560 1429.610 16.620 ;
        RECT 1299.110 16.420 1429.610 16.560 ;
        RECT 1299.110 16.360 1299.430 16.420 ;
        RECT 1429.290 16.360 1429.610 16.420 ;
      LAYER via ;
        RECT 1260.960 1322.640 1261.220 1322.900 ;
        RECT 1429.320 1315.160 1429.580 1315.420 ;
        RECT 1299.140 16.360 1299.400 16.620 ;
        RECT 1429.320 16.360 1429.580 16.620 ;
      LAYER met2 ;
        RECT 1259.530 1323.010 1259.810 1325.025 ;
        RECT 1259.530 1322.930 1261.160 1323.010 ;
        RECT 1259.530 1322.870 1261.220 1322.930 ;
        RECT 1259.530 1321.025 1259.810 1322.870 ;
        RECT 1260.960 1322.610 1261.220 1322.870 ;
        RECT 1429.320 1315.130 1429.580 1315.450 ;
        RECT 1429.380 16.650 1429.520 1315.130 ;
        RECT 1299.140 16.330 1299.400 16.650 ;
        RECT 1429.320 16.330 1429.580 16.650 ;
        RECT 1299.200 2.400 1299.340 16.330 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1317.050 176.700 1317.370 176.760 ;
        RECT 1418.710 176.700 1419.030 176.760 ;
        RECT 1317.050 176.560 1419.030 176.700 ;
        RECT 1317.050 176.500 1317.370 176.560 ;
        RECT 1418.710 176.500 1419.030 176.560 ;
      LAYER via ;
        RECT 1317.080 176.500 1317.340 176.760 ;
        RECT 1418.740 176.500 1419.000 176.760 ;
      LAYER met2 ;
        RECT 1418.730 482.955 1419.010 483.325 ;
        RECT 1418.800 176.790 1418.940 482.955 ;
        RECT 1317.080 176.470 1317.340 176.790 ;
        RECT 1418.740 176.470 1419.000 176.790 ;
        RECT 1317.140 2.400 1317.280 176.470 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
      LAYER via2 ;
        RECT 1418.730 483.000 1419.010 483.280 ;
      LAYER met3 ;
        RECT 1418.705 483.290 1419.035 483.305 ;
        RECT 1408.060 483.200 1419.035 483.290 ;
        RECT 1404.305 482.990 1419.035 483.200 ;
        RECT 1404.305 482.600 1408.305 482.990 ;
        RECT 1418.705 482.975 1419.035 482.990 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1264.150 1338.820 1264.470 1338.880 ;
        RECT 1421.930 1338.820 1422.250 1338.880 ;
        RECT 1264.150 1338.680 1422.250 1338.820 ;
        RECT 1264.150 1338.620 1264.470 1338.680 ;
        RECT 1421.930 1338.620 1422.250 1338.680 ;
        RECT 1334.990 30.160 1335.310 30.220 ;
        RECT 1421.930 30.160 1422.250 30.220 ;
        RECT 1334.990 30.020 1422.250 30.160 ;
        RECT 1334.990 29.960 1335.310 30.020 ;
        RECT 1421.930 29.960 1422.250 30.020 ;
      LAYER via ;
        RECT 1264.180 1338.620 1264.440 1338.880 ;
        RECT 1421.960 1338.620 1422.220 1338.880 ;
        RECT 1335.020 29.960 1335.280 30.220 ;
        RECT 1421.960 29.960 1422.220 30.220 ;
      LAYER met2 ;
        RECT 1264.180 1338.590 1264.440 1338.910 ;
        RECT 1421.960 1338.590 1422.220 1338.910 ;
        RECT 1264.240 1325.025 1264.380 1338.590 ;
        RECT 1264.130 1321.025 1264.410 1325.025 ;
        RECT 1422.020 30.250 1422.160 1338.590 ;
        RECT 1335.020 29.930 1335.280 30.250 ;
        RECT 1421.960 29.930 1422.220 30.250 ;
        RECT 1335.080 2.400 1335.220 29.930 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 692.370 17.240 692.690 17.300 ;
        RECT 696.510 17.240 696.830 17.300 ;
        RECT 692.370 17.100 696.830 17.240 ;
        RECT 692.370 17.040 692.690 17.100 ;
        RECT 696.510 17.040 696.830 17.100 ;
      LAYER via ;
        RECT 692.400 17.040 692.660 17.300 ;
        RECT 696.540 17.040 696.800 17.300 ;
      LAYER met2 ;
        RECT 1415.970 1206.475 1416.250 1206.845 ;
        RECT 1416.040 263.005 1416.180 1206.475 ;
        RECT 1415.970 262.635 1416.250 263.005 ;
        RECT 696.530 149.075 696.810 149.445 ;
        RECT 696.600 17.330 696.740 149.075 ;
        RECT 692.400 17.010 692.660 17.330 ;
        RECT 696.540 17.010 696.800 17.330 ;
        RECT 692.460 2.400 692.600 17.010 ;
        RECT 692.250 -4.800 692.810 2.400 ;
      LAYER via2 ;
        RECT 1415.970 1206.520 1416.250 1206.800 ;
        RECT 1415.970 262.680 1416.250 262.960 ;
        RECT 696.530 149.120 696.810 149.400 ;
      LAYER met3 ;
        RECT 1415.945 1206.810 1416.275 1206.825 ;
        RECT 1408.060 1206.720 1416.275 1206.810 ;
        RECT 1404.305 1206.510 1416.275 1206.720 ;
        RECT 1404.305 1206.120 1408.305 1206.510 ;
        RECT 1415.945 1206.495 1416.275 1206.510 ;
        RECT 1415.945 262.980 1416.275 262.985 ;
        RECT 1415.945 262.970 1416.530 262.980 ;
        RECT 1415.720 262.670 1416.530 262.970 ;
        RECT 1415.945 262.660 1416.530 262.670 ;
        RECT 1415.945 262.655 1416.275 262.660 ;
        RECT 696.505 149.410 696.835 149.425 ;
        RECT 1416.150 149.410 1416.530 149.420 ;
        RECT 696.505 149.110 1416.530 149.410 ;
        RECT 696.505 149.095 696.835 149.110 ;
        RECT 1416.150 149.100 1416.530 149.110 ;
      LAYER via3 ;
        RECT 1416.180 262.660 1416.500 262.980 ;
        RECT 1416.180 149.100 1416.500 149.420 ;
      LAYER met4 ;
        RECT 1416.175 262.655 1416.505 262.985 ;
        RECT 1416.190 149.425 1416.490 262.655 ;
        RECT 1416.175 149.095 1416.505 149.425 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 895.690 162.760 896.010 162.820 ;
        RECT 1352.470 162.760 1352.790 162.820 ;
        RECT 895.690 162.620 1352.790 162.760 ;
        RECT 895.690 162.560 896.010 162.620 ;
        RECT 1352.470 162.560 1352.790 162.620 ;
      LAYER via ;
        RECT 895.720 162.560 895.980 162.820 ;
        RECT 1352.500 162.560 1352.760 162.820 ;
      LAYER met2 ;
        RECT 896.130 216.650 896.410 220.000 ;
        RECT 895.780 216.510 896.410 216.650 ;
        RECT 895.780 162.850 895.920 216.510 ;
        RECT 896.130 216.000 896.410 216.510 ;
        RECT 895.720 162.530 895.980 162.850 ;
        RECT 1352.500 162.530 1352.760 162.850 ;
        RECT 1352.560 2.400 1352.700 162.530 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 713.070 200.500 713.390 200.560 ;
        RECT 717.210 200.500 717.530 200.560 ;
        RECT 713.070 200.360 717.530 200.500 ;
        RECT 713.070 200.300 713.390 200.360 ;
        RECT 717.210 200.300 717.530 200.360 ;
        RECT 717.210 25.060 717.530 25.120 ;
        RECT 1370.410 25.060 1370.730 25.120 ;
        RECT 717.210 24.920 1370.730 25.060 ;
        RECT 717.210 24.860 717.530 24.920 ;
        RECT 1370.410 24.860 1370.730 24.920 ;
      LAYER via ;
        RECT 713.100 200.300 713.360 200.560 ;
        RECT 717.240 200.300 717.500 200.560 ;
        RECT 717.240 24.860 717.500 25.120 ;
        RECT 1370.440 24.860 1370.700 25.120 ;
      LAYER met2 ;
        RECT 713.050 216.000 713.330 220.000 ;
        RECT 713.160 200.590 713.300 216.000 ;
        RECT 713.100 200.270 713.360 200.590 ;
        RECT 717.240 200.270 717.500 200.590 ;
        RECT 717.300 25.150 717.440 200.270 ;
        RECT 717.240 24.830 717.500 25.150 ;
        RECT 1370.440 24.830 1370.700 25.150 ;
        RECT 1370.500 2.400 1370.640 24.830 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 824.390 1348.680 824.710 1348.740 ;
        RECT 1442.630 1348.680 1442.950 1348.740 ;
        RECT 824.390 1348.540 1442.950 1348.680 ;
        RECT 824.390 1348.480 824.710 1348.540 ;
        RECT 1442.630 1348.480 1442.950 1348.540 ;
        RECT 1388.350 29.820 1388.670 29.880 ;
        RECT 1442.630 29.820 1442.950 29.880 ;
        RECT 1388.350 29.680 1442.950 29.820 ;
        RECT 1388.350 29.620 1388.670 29.680 ;
        RECT 1442.630 29.620 1442.950 29.680 ;
      LAYER via ;
        RECT 824.420 1348.480 824.680 1348.740 ;
        RECT 1442.660 1348.480 1442.920 1348.740 ;
        RECT 1388.380 29.620 1388.640 29.880 ;
        RECT 1442.660 29.620 1442.920 29.880 ;
      LAYER met2 ;
        RECT 824.420 1348.450 824.680 1348.770 ;
        RECT 1442.660 1348.450 1442.920 1348.770 ;
        RECT 824.480 1325.025 824.620 1348.450 ;
        RECT 824.370 1321.025 824.650 1325.025 ;
        RECT 1442.720 29.910 1442.860 1348.450 ;
        RECT 1388.380 29.590 1388.640 29.910 ;
        RECT 1442.660 29.590 1442.920 29.910 ;
        RECT 1388.440 2.400 1388.580 29.590 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 295.850 120.940 296.170 121.000 ;
        RECT 1400.770 120.940 1401.090 121.000 ;
        RECT 295.850 120.800 1401.090 120.940 ;
        RECT 295.850 120.740 296.170 120.800 ;
        RECT 1400.770 120.740 1401.090 120.800 ;
        RECT 1400.770 2.960 1401.090 3.020 ;
        RECT 1406.290 2.960 1406.610 3.020 ;
        RECT 1400.770 2.820 1406.610 2.960 ;
        RECT 1400.770 2.760 1401.090 2.820 ;
        RECT 1406.290 2.760 1406.610 2.820 ;
      LAYER via ;
        RECT 295.880 120.740 296.140 121.000 ;
        RECT 1400.800 120.740 1401.060 121.000 ;
        RECT 1400.800 2.760 1401.060 3.020 ;
        RECT 1406.320 2.760 1406.580 3.020 ;
      LAYER met2 ;
        RECT 295.870 1169.755 296.150 1170.125 ;
        RECT 295.940 121.030 296.080 1169.755 ;
        RECT 295.880 120.710 296.140 121.030 ;
        RECT 1400.800 120.710 1401.060 121.030 ;
        RECT 1400.860 3.050 1401.000 120.710 ;
        RECT 1400.800 2.730 1401.060 3.050 ;
        RECT 1406.320 2.730 1406.580 3.050 ;
        RECT 1406.380 2.400 1406.520 2.730 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
      LAYER via2 ;
        RECT 295.870 1169.800 296.150 1170.080 ;
      LAYER met3 ;
        RECT 295.845 1170.090 296.175 1170.105 ;
        RECT 295.845 1170.000 310.500 1170.090 ;
        RECT 295.845 1169.790 314.000 1170.000 ;
        RECT 295.845 1169.775 296.175 1169.790 ;
        RECT 310.000 1169.400 314.000 1169.790 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1155.590 1328.960 1155.910 1329.020 ;
        RECT 1421.470 1328.960 1421.790 1329.020 ;
        RECT 1155.590 1328.820 1421.790 1328.960 ;
        RECT 1155.590 1328.760 1155.910 1328.820 ;
        RECT 1421.470 1328.760 1421.790 1328.820 ;
      LAYER via ;
        RECT 1155.620 1328.760 1155.880 1329.020 ;
        RECT 1421.500 1328.760 1421.760 1329.020 ;
      LAYER met2 ;
        RECT 1155.620 1328.730 1155.880 1329.050 ;
        RECT 1421.500 1328.730 1421.760 1329.050 ;
        RECT 1155.680 1325.025 1155.820 1328.730 ;
        RECT 1155.570 1321.025 1155.850 1325.025 ;
        RECT 1421.560 17.410 1421.700 1328.730 ;
        RECT 1421.560 17.270 1424.000 17.410 ;
        RECT 1423.860 2.400 1424.000 17.270 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1344.650 1324.880 1344.970 1324.940 ;
        RECT 1435.270 1324.880 1435.590 1324.940 ;
        RECT 1344.650 1324.740 1435.590 1324.880 ;
        RECT 1344.650 1324.680 1344.970 1324.740 ;
        RECT 1435.270 1324.680 1435.590 1324.740 ;
        RECT 1435.270 16.900 1435.590 16.960 ;
        RECT 1441.710 16.900 1442.030 16.960 ;
        RECT 1435.270 16.760 1442.030 16.900 ;
        RECT 1435.270 16.700 1435.590 16.760 ;
        RECT 1441.710 16.700 1442.030 16.760 ;
      LAYER via ;
        RECT 1344.680 1324.680 1344.940 1324.940 ;
        RECT 1435.300 1324.680 1435.560 1324.940 ;
        RECT 1435.300 16.700 1435.560 16.960 ;
        RECT 1441.740 16.700 1442.000 16.960 ;
      LAYER met2 ;
        RECT 1343.430 1325.025 1344.880 1325.050 ;
        RECT 1343.250 1324.970 1344.880 1325.025 ;
        RECT 1343.250 1324.910 1344.940 1324.970 ;
        RECT 1343.250 1321.025 1343.530 1324.910 ;
        RECT 1344.680 1324.650 1344.940 1324.910 ;
        RECT 1435.300 1324.650 1435.560 1324.970 ;
        RECT 1435.360 16.990 1435.500 1324.650 ;
        RECT 1435.300 16.670 1435.560 16.990 ;
        RECT 1441.740 16.670 1442.000 16.990 ;
        RECT 1441.800 2.400 1441.940 16.670 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1346.030 200.500 1346.350 200.560 ;
        RECT 1352.010 200.500 1352.330 200.560 ;
        RECT 1346.030 200.360 1352.330 200.500 ;
        RECT 1346.030 200.300 1346.350 200.360 ;
        RECT 1352.010 200.300 1352.330 200.360 ;
        RECT 1352.010 80.480 1352.330 80.540 ;
        RECT 1455.970 80.480 1456.290 80.540 ;
        RECT 1352.010 80.340 1456.290 80.480 ;
        RECT 1352.010 80.280 1352.330 80.340 ;
        RECT 1455.970 80.280 1456.290 80.340 ;
      LAYER via ;
        RECT 1346.060 200.300 1346.320 200.560 ;
        RECT 1352.040 200.300 1352.300 200.560 ;
        RECT 1352.040 80.280 1352.300 80.540 ;
        RECT 1456.000 80.280 1456.260 80.540 ;
      LAYER met2 ;
        RECT 1346.010 216.000 1346.290 220.000 ;
        RECT 1346.120 200.590 1346.260 216.000 ;
        RECT 1346.060 200.270 1346.320 200.590 ;
        RECT 1352.040 200.270 1352.300 200.590 ;
        RECT 1352.100 80.570 1352.240 200.270 ;
        RECT 1352.040 80.250 1352.300 80.570 ;
        RECT 1456.000 80.250 1456.260 80.570 ;
        RECT 1456.060 16.730 1456.200 80.250 ;
        RECT 1456.060 16.590 1459.880 16.730 ;
        RECT 1459.740 2.400 1459.880 16.590 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 292.630 655.760 292.950 655.820 ;
        RECT 296.770 655.760 297.090 655.820 ;
        RECT 292.630 655.620 297.090 655.760 ;
        RECT 292.630 655.560 292.950 655.620 ;
        RECT 296.770 655.560 297.090 655.620 ;
        RECT 292.630 155.960 292.950 156.020 ;
        RECT 1476.670 155.960 1476.990 156.020 ;
        RECT 292.630 155.820 1476.990 155.960 ;
        RECT 292.630 155.760 292.950 155.820 ;
        RECT 1476.670 155.760 1476.990 155.820 ;
      LAYER via ;
        RECT 292.660 655.560 292.920 655.820 ;
        RECT 296.800 655.560 297.060 655.820 ;
        RECT 292.660 155.760 292.920 156.020 ;
        RECT 1476.700 155.760 1476.960 156.020 ;
      LAYER met2 ;
        RECT 296.790 658.395 297.070 658.765 ;
        RECT 296.860 655.850 297.000 658.395 ;
        RECT 292.660 655.530 292.920 655.850 ;
        RECT 296.800 655.530 297.060 655.850 ;
        RECT 292.720 156.050 292.860 655.530 ;
        RECT 292.660 155.730 292.920 156.050 ;
        RECT 1476.700 155.730 1476.960 156.050 ;
        RECT 1476.760 16.730 1476.900 155.730 ;
        RECT 1476.760 16.590 1477.820 16.730 ;
        RECT 1477.680 2.400 1477.820 16.590 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
      LAYER via2 ;
        RECT 296.790 658.440 297.070 658.720 ;
      LAYER met3 ;
        RECT 296.765 658.730 297.095 658.745 ;
        RECT 296.765 658.640 310.500 658.730 ;
        RECT 296.765 658.430 314.000 658.640 ;
        RECT 296.765 658.415 297.095 658.430 ;
        RECT 310.000 658.040 314.000 658.430 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1105.910 1327.260 1106.230 1327.320 ;
        RECT 1490.470 1327.260 1490.790 1327.320 ;
        RECT 1105.910 1327.120 1490.790 1327.260 ;
        RECT 1105.910 1327.060 1106.230 1327.120 ;
        RECT 1490.470 1327.060 1490.790 1327.120 ;
      LAYER via ;
        RECT 1105.940 1327.060 1106.200 1327.320 ;
        RECT 1490.500 1327.060 1490.760 1327.320 ;
      LAYER met2 ;
        RECT 1105.940 1327.030 1106.200 1327.350 ;
        RECT 1490.500 1327.030 1490.760 1327.350 ;
        RECT 1106.000 1325.025 1106.140 1327.030 ;
        RECT 1105.890 1321.025 1106.170 1325.025 ;
        RECT 1490.560 17.410 1490.700 1327.030 ;
        RECT 1490.560 17.270 1495.760 17.410 ;
        RECT 1495.620 2.400 1495.760 17.270 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1242.260 1421.330 1242.320 ;
        RECT 1511.170 1242.260 1511.490 1242.320 ;
        RECT 1421.010 1242.120 1511.490 1242.260 ;
        RECT 1421.010 1242.060 1421.330 1242.120 ;
        RECT 1511.170 1242.060 1511.490 1242.120 ;
      LAYER via ;
        RECT 1421.040 1242.060 1421.300 1242.320 ;
        RECT 1511.200 1242.060 1511.460 1242.320 ;
      LAYER met2 ;
        RECT 1421.030 1243.195 1421.310 1243.565 ;
        RECT 1421.100 1242.350 1421.240 1243.195 ;
        RECT 1421.040 1242.030 1421.300 1242.350 ;
        RECT 1511.200 1242.030 1511.460 1242.350 ;
        RECT 1511.260 17.410 1511.400 1242.030 ;
        RECT 1511.260 17.270 1513.240 17.410 ;
        RECT 1513.100 2.400 1513.240 17.270 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1243.240 1421.310 1243.520 ;
      LAYER met3 ;
        RECT 1421.005 1243.530 1421.335 1243.545 ;
        RECT 1408.060 1243.440 1421.335 1243.530 ;
        RECT 1404.305 1243.230 1421.335 1243.440 ;
        RECT 1404.305 1242.840 1408.305 1243.230 ;
        RECT 1421.005 1243.215 1421.335 1243.230 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 472.565 15.385 472.735 17.255 ;
        RECT 520.865 15.385 521.035 17.595 ;
        RECT 641.845 16.065 642.015 17.255 ;
      LAYER mcon ;
        RECT 520.865 17.425 521.035 17.595 ;
        RECT 472.565 17.085 472.735 17.255 ;
        RECT 641.845 17.085 642.015 17.255 ;
      LAYER met1 ;
        RECT 275.610 1332.360 275.930 1332.420 ;
        RECT 334.950 1332.360 335.270 1332.420 ;
        RECT 275.610 1332.220 335.270 1332.360 ;
        RECT 275.610 1332.160 275.930 1332.220 ;
        RECT 334.950 1332.160 335.270 1332.220 ;
        RECT 520.805 17.580 521.095 17.625 ;
        RECT 520.805 17.440 569.780 17.580 ;
        RECT 520.805 17.395 521.095 17.440 ;
        RECT 275.610 17.240 275.930 17.300 ;
        RECT 472.505 17.240 472.795 17.285 ;
        RECT 275.610 17.100 472.795 17.240 ;
        RECT 275.610 17.040 275.930 17.100 ;
        RECT 472.505 17.055 472.795 17.100 ;
        RECT 569.640 16.900 569.780 17.440 ;
        RECT 641.785 17.240 642.075 17.285 ;
        RECT 613.340 17.100 642.075 17.240 ;
        RECT 613.340 16.900 613.480 17.100 ;
        RECT 641.785 17.055 642.075 17.100 ;
        RECT 569.640 16.760 613.480 16.900 ;
        RECT 641.785 16.220 642.075 16.265 ;
        RECT 710.310 16.220 710.630 16.280 ;
        RECT 641.785 16.080 710.630 16.220 ;
        RECT 641.785 16.035 642.075 16.080 ;
        RECT 710.310 16.020 710.630 16.080 ;
        RECT 472.505 15.540 472.795 15.585 ;
        RECT 520.805 15.540 521.095 15.585 ;
        RECT 472.505 15.400 521.095 15.540 ;
        RECT 472.505 15.355 472.795 15.400 ;
        RECT 520.805 15.355 521.095 15.400 ;
      LAYER via ;
        RECT 275.640 1332.160 275.900 1332.420 ;
        RECT 334.980 1332.160 335.240 1332.420 ;
        RECT 275.640 17.040 275.900 17.300 ;
        RECT 710.340 16.020 710.600 16.280 ;
      LAYER met2 ;
        RECT 275.640 1332.130 275.900 1332.450 ;
        RECT 334.980 1332.130 335.240 1332.450 ;
        RECT 275.700 17.330 275.840 1332.130 ;
        RECT 335.040 1325.025 335.180 1332.130 ;
        RECT 334.930 1321.025 335.210 1325.025 ;
        RECT 275.640 17.010 275.900 17.330 ;
        RECT 710.340 15.990 710.600 16.310 ;
        RECT 710.400 2.400 710.540 15.990 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1217.230 200.500 1217.550 200.560 ;
        RECT 1220.910 200.500 1221.230 200.560 ;
        RECT 1217.230 200.360 1221.230 200.500 ;
        RECT 1217.230 200.300 1217.550 200.360 ;
        RECT 1220.910 200.300 1221.230 200.360 ;
        RECT 1220.910 30.500 1221.230 30.560 ;
        RECT 1530.950 30.500 1531.270 30.560 ;
        RECT 1220.910 30.360 1531.270 30.500 ;
        RECT 1220.910 30.300 1221.230 30.360 ;
        RECT 1530.950 30.300 1531.270 30.360 ;
      LAYER via ;
        RECT 1217.260 200.300 1217.520 200.560 ;
        RECT 1220.940 200.300 1221.200 200.560 ;
        RECT 1220.940 30.300 1221.200 30.560 ;
        RECT 1530.980 30.300 1531.240 30.560 ;
      LAYER met2 ;
        RECT 1217.210 216.000 1217.490 220.000 ;
        RECT 1217.320 200.590 1217.460 216.000 ;
        RECT 1217.260 200.270 1217.520 200.590 ;
        RECT 1220.940 200.270 1221.200 200.590 ;
        RECT 1221.000 30.590 1221.140 200.270 ;
        RECT 1220.940 30.270 1221.200 30.590 ;
        RECT 1530.980 30.270 1531.240 30.590 ;
        RECT 1531.040 2.400 1531.180 30.270 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 296.310 80.140 296.630 80.200 ;
        RECT 1545.670 80.140 1545.990 80.200 ;
        RECT 296.310 80.000 1545.990 80.140 ;
        RECT 296.310 79.940 296.630 80.000 ;
        RECT 1545.670 79.940 1545.990 80.000 ;
      LAYER via ;
        RECT 296.340 79.940 296.600 80.200 ;
        RECT 1545.700 79.940 1545.960 80.200 ;
      LAYER met2 ;
        RECT 296.330 1199.675 296.610 1200.045 ;
        RECT 296.400 80.230 296.540 1199.675 ;
        RECT 296.340 79.910 296.600 80.230 ;
        RECT 1545.700 79.910 1545.960 80.230 ;
        RECT 1545.760 17.410 1545.900 79.910 ;
        RECT 1545.760 17.270 1549.120 17.410 ;
        RECT 1548.980 2.400 1549.120 17.270 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
      LAYER via2 ;
        RECT 296.330 1199.720 296.610 1200.000 ;
      LAYER met3 ;
        RECT 296.305 1200.010 296.635 1200.025 ;
        RECT 296.305 1199.920 310.500 1200.010 ;
        RECT 296.305 1199.710 314.000 1199.920 ;
        RECT 296.305 1199.695 296.635 1199.710 ;
        RECT 310.000 1199.320 314.000 1199.710 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1152.830 200.500 1153.150 200.560 ;
        RECT 1158.810 200.500 1159.130 200.560 ;
        RECT 1152.830 200.360 1159.130 200.500 ;
        RECT 1152.830 200.300 1153.150 200.360 ;
        RECT 1158.810 200.300 1159.130 200.360 ;
        RECT 1158.810 143.040 1159.130 143.100 ;
        RECT 1566.830 143.040 1567.150 143.100 ;
        RECT 1158.810 142.900 1567.150 143.040 ;
        RECT 1158.810 142.840 1159.130 142.900 ;
        RECT 1566.830 142.840 1567.150 142.900 ;
      LAYER via ;
        RECT 1152.860 200.300 1153.120 200.560 ;
        RECT 1158.840 200.300 1159.100 200.560 ;
        RECT 1158.840 142.840 1159.100 143.100 ;
        RECT 1566.860 142.840 1567.120 143.100 ;
      LAYER met2 ;
        RECT 1152.810 216.000 1153.090 220.000 ;
        RECT 1152.920 200.590 1153.060 216.000 ;
        RECT 1152.860 200.270 1153.120 200.590 ;
        RECT 1158.840 200.270 1159.100 200.590 ;
        RECT 1158.900 143.130 1159.040 200.270 ;
        RECT 1158.840 142.810 1159.100 143.130 ;
        RECT 1566.860 142.810 1567.120 143.130 ;
        RECT 1566.920 2.400 1567.060 142.810 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1416.870 800.600 1417.190 800.660 ;
        RECT 1580.170 800.600 1580.490 800.660 ;
        RECT 1416.870 800.460 1580.490 800.600 ;
        RECT 1416.870 800.400 1417.190 800.460 ;
        RECT 1580.170 800.400 1580.490 800.460 ;
        RECT 1580.170 2.960 1580.490 3.020 ;
        RECT 1584.770 2.960 1585.090 3.020 ;
        RECT 1580.170 2.820 1585.090 2.960 ;
        RECT 1580.170 2.760 1580.490 2.820 ;
        RECT 1584.770 2.760 1585.090 2.820 ;
      LAYER via ;
        RECT 1416.900 800.400 1417.160 800.660 ;
        RECT 1580.200 800.400 1580.460 800.660 ;
        RECT 1580.200 2.760 1580.460 3.020 ;
        RECT 1584.800 2.760 1585.060 3.020 ;
      LAYER met2 ;
        RECT 1416.890 805.275 1417.170 805.645 ;
        RECT 1416.960 800.690 1417.100 805.275 ;
        RECT 1416.900 800.370 1417.160 800.690 ;
        RECT 1580.200 800.370 1580.460 800.690 ;
        RECT 1580.260 3.050 1580.400 800.370 ;
        RECT 1580.200 2.730 1580.460 3.050 ;
        RECT 1584.800 2.730 1585.060 3.050 ;
        RECT 1584.860 2.400 1585.000 2.730 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
      LAYER via2 ;
        RECT 1416.890 805.320 1417.170 805.600 ;
      LAYER met3 ;
        RECT 1416.865 805.610 1417.195 805.625 ;
        RECT 1408.060 805.520 1417.195 805.610 ;
        RECT 1404.305 805.310 1417.195 805.520 ;
        RECT 1404.305 804.920 1408.305 805.310 ;
        RECT 1416.865 805.295 1417.195 805.310 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1269.210 107.680 1269.530 107.740 ;
        RECT 1600.870 107.680 1601.190 107.740 ;
        RECT 1269.210 107.540 1601.190 107.680 ;
        RECT 1269.210 107.480 1269.530 107.540 ;
        RECT 1600.870 107.480 1601.190 107.540 ;
      LAYER via ;
        RECT 1269.240 107.480 1269.500 107.740 ;
        RECT 1600.900 107.480 1601.160 107.740 ;
      LAYER met2 ;
        RECT 1266.890 216.650 1267.170 220.000 ;
        RECT 1266.890 216.510 1269.440 216.650 ;
        RECT 1266.890 216.000 1267.170 216.510 ;
        RECT 1269.300 107.770 1269.440 216.510 ;
        RECT 1269.240 107.450 1269.500 107.770 ;
        RECT 1600.900 107.450 1601.160 107.770 ;
        RECT 1600.960 3.130 1601.100 107.450 ;
        RECT 1600.960 2.990 1602.480 3.130 ;
        RECT 1602.340 2.400 1602.480 2.990 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 436.150 204.240 436.470 204.300 ;
        RECT 1614.670 204.240 1614.990 204.300 ;
        RECT 436.150 204.100 1614.990 204.240 ;
        RECT 436.150 204.040 436.470 204.100 ;
        RECT 1614.670 204.040 1614.990 204.100 ;
        RECT 1614.670 2.960 1614.990 3.020 ;
        RECT 1620.190 2.960 1620.510 3.020 ;
        RECT 1614.670 2.820 1620.510 2.960 ;
        RECT 1614.670 2.760 1614.990 2.820 ;
        RECT 1620.190 2.760 1620.510 2.820 ;
      LAYER via ;
        RECT 436.180 204.040 436.440 204.300 ;
        RECT 1614.700 204.040 1614.960 204.300 ;
        RECT 1614.700 2.760 1614.960 3.020 ;
        RECT 1620.220 2.760 1620.480 3.020 ;
      LAYER met2 ;
        RECT 436.130 216.000 436.410 220.000 ;
        RECT 436.240 204.330 436.380 216.000 ;
        RECT 436.180 204.010 436.440 204.330 ;
        RECT 1614.700 204.010 1614.960 204.330 ;
        RECT 1614.760 3.050 1614.900 204.010 ;
        RECT 1614.700 2.730 1614.960 3.050 ;
        RECT 1620.220 2.730 1620.480 3.050 ;
        RECT 1620.280 2.400 1620.420 2.730 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 1326.580 483.390 1326.640 ;
        RECT 1635.370 1326.580 1635.690 1326.640 ;
        RECT 483.070 1326.440 1635.690 1326.580 ;
        RECT 483.070 1326.380 483.390 1326.440 ;
        RECT 1635.370 1326.380 1635.690 1326.440 ;
      LAYER via ;
        RECT 483.100 1326.380 483.360 1326.640 ;
        RECT 1635.400 1326.380 1635.660 1326.640 ;
      LAYER met2 ;
        RECT 483.100 1326.350 483.360 1326.670 ;
        RECT 1635.400 1326.350 1635.660 1326.670 ;
        RECT 483.160 1325.025 483.300 1326.350 ;
        RECT 483.050 1321.025 483.330 1325.025 ;
        RECT 1635.460 17.410 1635.600 1326.350 ;
        RECT 1635.460 17.270 1638.360 17.410 ;
        RECT 1638.220 2.400 1638.360 17.270 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1062.740 1421.330 1062.800 ;
        RECT 1656.070 1062.740 1656.390 1062.800 ;
        RECT 1421.010 1062.600 1656.390 1062.740 ;
        RECT 1421.010 1062.540 1421.330 1062.600 ;
        RECT 1656.070 1062.540 1656.390 1062.600 ;
      LAYER via ;
        RECT 1421.040 1062.540 1421.300 1062.800 ;
        RECT 1656.100 1062.540 1656.360 1062.800 ;
      LAYER met2 ;
        RECT 1421.030 1067.755 1421.310 1068.125 ;
        RECT 1421.100 1062.830 1421.240 1067.755 ;
        RECT 1421.040 1062.510 1421.300 1062.830 ;
        RECT 1656.100 1062.510 1656.360 1062.830 ;
        RECT 1656.160 2.400 1656.300 1062.510 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1067.800 1421.310 1068.080 ;
      LAYER met3 ;
        RECT 1421.005 1068.090 1421.335 1068.105 ;
        RECT 1408.060 1068.000 1421.335 1068.090 ;
        RECT 1404.305 1067.790 1421.335 1068.000 ;
        RECT 1404.305 1067.400 1408.305 1067.790 ;
        RECT 1421.005 1067.775 1421.335 1067.790 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 301.370 217.500 301.690 217.560 ;
        RECT 1669.870 217.500 1670.190 217.560 ;
        RECT 301.370 217.360 1670.190 217.500 ;
        RECT 301.370 217.300 301.690 217.360 ;
        RECT 1669.870 217.300 1670.190 217.360 ;
      LAYER via ;
        RECT 301.400 217.300 301.660 217.560 ;
        RECT 1669.900 217.300 1670.160 217.560 ;
      LAYER met2 ;
        RECT 301.390 526.475 301.670 526.845 ;
        RECT 301.460 217.590 301.600 526.475 ;
        RECT 301.400 217.270 301.660 217.590 ;
        RECT 1669.900 217.270 1670.160 217.590 ;
        RECT 1669.960 17.410 1670.100 217.270 ;
        RECT 1669.960 17.270 1673.780 17.410 ;
        RECT 1673.640 2.400 1673.780 17.270 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
      LAYER via2 ;
        RECT 301.390 526.520 301.670 526.800 ;
      LAYER met3 ;
        RECT 301.365 526.810 301.695 526.825 ;
        RECT 301.365 526.720 310.500 526.810 ;
        RECT 301.365 526.510 314.000 526.720 ;
        RECT 301.365 526.495 301.695 526.510 ;
        RECT 310.000 526.120 314.000 526.510 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1350.630 206.620 1350.950 206.680 ;
        RECT 1690.570 206.620 1690.890 206.680 ;
        RECT 1350.630 206.480 1690.890 206.620 ;
        RECT 1350.630 206.420 1350.950 206.480 ;
        RECT 1690.570 206.420 1690.890 206.480 ;
      LAYER via ;
        RECT 1350.660 206.420 1350.920 206.680 ;
        RECT 1690.600 206.420 1690.860 206.680 ;
      LAYER met2 ;
        RECT 1350.610 216.000 1350.890 220.000 ;
        RECT 1350.720 206.710 1350.860 216.000 ;
        RECT 1350.660 206.390 1350.920 206.710 ;
        RECT 1690.600 206.390 1690.860 206.710 ;
        RECT 1690.660 17.410 1690.800 206.390 ;
        RECT 1690.660 17.270 1691.720 17.410 ;
        RECT 1691.580 2.400 1691.720 17.270 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 302.290 219.200 302.610 219.260 ;
        RECT 720.890 219.200 721.210 219.260 ;
        RECT 302.290 219.060 721.210 219.200 ;
        RECT 302.290 219.000 302.610 219.060 ;
        RECT 720.890 219.000 721.210 219.060 ;
        RECT 720.890 17.240 721.210 17.300 ;
        RECT 728.250 17.240 728.570 17.300 ;
        RECT 720.890 17.100 728.570 17.240 ;
        RECT 720.890 17.040 721.210 17.100 ;
        RECT 728.250 17.040 728.570 17.100 ;
      LAYER via ;
        RECT 302.320 219.000 302.580 219.260 ;
        RECT 720.920 219.000 721.180 219.260 ;
        RECT 720.920 17.040 721.180 17.300 ;
        RECT 728.280 17.040 728.540 17.300 ;
      LAYER met2 ;
        RECT 302.310 247.675 302.590 248.045 ;
        RECT 302.380 219.290 302.520 247.675 ;
        RECT 302.320 218.970 302.580 219.290 ;
        RECT 720.920 218.970 721.180 219.290 ;
        RECT 720.980 17.330 721.120 218.970 ;
        RECT 720.920 17.010 721.180 17.330 ;
        RECT 728.280 17.010 728.540 17.330 ;
        RECT 728.340 2.400 728.480 17.010 ;
        RECT 728.130 -4.800 728.690 2.400 ;
      LAYER via2 ;
        RECT 302.310 247.720 302.590 248.000 ;
      LAYER met3 ;
        RECT 310.000 248.690 314.000 249.280 ;
        RECT 302.990 248.680 314.000 248.690 ;
        RECT 302.990 248.390 310.650 248.680 ;
        RECT 302.285 248.010 302.615 248.025 ;
        RECT 302.990 248.010 303.290 248.390 ;
        RECT 302.285 247.710 303.290 248.010 ;
        RECT 302.285 247.695 302.615 247.710 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 294.470 176.360 294.790 176.420 ;
        RECT 1704.370 176.360 1704.690 176.420 ;
        RECT 294.470 176.220 1704.690 176.360 ;
        RECT 294.470 176.160 294.790 176.220 ;
        RECT 1704.370 176.160 1704.690 176.220 ;
      LAYER via ;
        RECT 294.500 176.160 294.760 176.420 ;
        RECT 1704.400 176.160 1704.660 176.420 ;
      LAYER met2 ;
        RECT 294.490 935.835 294.770 936.205 ;
        RECT 294.560 176.450 294.700 935.835 ;
        RECT 294.500 176.130 294.760 176.450 ;
        RECT 1704.400 176.130 1704.660 176.450 ;
        RECT 1704.460 17.410 1704.600 176.130 ;
        RECT 1704.460 17.270 1709.660 17.410 ;
        RECT 1709.520 2.400 1709.660 17.270 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
      LAYER via2 ;
        RECT 294.490 935.880 294.770 936.160 ;
      LAYER met3 ;
        RECT 294.465 936.170 294.795 936.185 ;
        RECT 294.465 936.080 310.500 936.170 ;
        RECT 294.465 935.870 314.000 936.080 ;
        RECT 294.465 935.855 294.795 935.870 ;
        RECT 310.000 935.480 314.000 935.870 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1378.230 1327.940 1378.550 1328.000 ;
        RECT 1725.070 1327.940 1725.390 1328.000 ;
        RECT 1378.230 1327.800 1725.390 1327.940 ;
        RECT 1378.230 1327.740 1378.550 1327.800 ;
        RECT 1725.070 1327.740 1725.390 1327.800 ;
      LAYER via ;
        RECT 1378.260 1327.740 1378.520 1328.000 ;
        RECT 1725.100 1327.740 1725.360 1328.000 ;
      LAYER met2 ;
        RECT 1378.260 1327.710 1378.520 1328.030 ;
        RECT 1725.100 1327.710 1725.360 1328.030 ;
        RECT 1378.320 1325.025 1378.460 1327.710 ;
        RECT 1378.210 1321.025 1378.490 1325.025 ;
        RECT 1725.160 17.410 1725.300 1327.710 ;
        RECT 1725.160 17.270 1727.600 17.410 ;
        RECT 1727.460 2.400 1727.600 17.270 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 344.150 1325.560 344.470 1325.620 ;
        RECT 1738.870 1325.560 1739.190 1325.620 ;
        RECT 344.150 1325.420 1739.190 1325.560 ;
        RECT 344.150 1325.360 344.470 1325.420 ;
        RECT 1738.870 1325.360 1739.190 1325.420 ;
        RECT 1738.870 16.900 1739.190 16.960 ;
        RECT 1745.310 16.900 1745.630 16.960 ;
        RECT 1738.870 16.760 1745.630 16.900 ;
        RECT 1738.870 16.700 1739.190 16.760 ;
        RECT 1745.310 16.700 1745.630 16.760 ;
      LAYER via ;
        RECT 344.180 1325.360 344.440 1325.620 ;
        RECT 1738.900 1325.360 1739.160 1325.620 ;
        RECT 1738.900 16.700 1739.160 16.960 ;
        RECT 1745.340 16.700 1745.600 16.960 ;
      LAYER met2 ;
        RECT 344.180 1325.330 344.440 1325.650 ;
        RECT 1738.900 1325.330 1739.160 1325.650 ;
        RECT 344.240 1325.025 344.380 1325.330 ;
        RECT 344.130 1321.025 344.410 1325.025 ;
        RECT 1738.960 16.990 1739.100 1325.330 ;
        RECT 1738.900 16.670 1739.160 16.990 ;
        RECT 1745.340 16.670 1745.600 16.990 ;
        RECT 1745.400 2.400 1745.540 16.670 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 611.870 1332.020 612.190 1332.080 ;
        RECT 641.770 1332.020 642.090 1332.080 ;
        RECT 611.870 1331.880 642.090 1332.020 ;
        RECT 611.870 1331.820 612.190 1331.880 ;
        RECT 641.770 1331.820 642.090 1331.880 ;
        RECT 641.770 1328.280 642.090 1328.340 ;
        RECT 1759.570 1328.280 1759.890 1328.340 ;
        RECT 641.770 1328.140 1759.890 1328.280 ;
        RECT 641.770 1328.080 642.090 1328.140 ;
        RECT 1759.570 1328.080 1759.890 1328.140 ;
      LAYER via ;
        RECT 611.900 1331.820 612.160 1332.080 ;
        RECT 641.800 1331.820 642.060 1332.080 ;
        RECT 641.800 1328.080 642.060 1328.340 ;
        RECT 1759.600 1328.080 1759.860 1328.340 ;
      LAYER met2 ;
        RECT 611.900 1331.790 612.160 1332.110 ;
        RECT 641.800 1331.790 642.060 1332.110 ;
        RECT 611.960 1325.025 612.100 1331.790 ;
        RECT 641.860 1328.370 642.000 1331.790 ;
        RECT 641.800 1328.050 642.060 1328.370 ;
        RECT 1759.600 1328.050 1759.860 1328.370 ;
        RECT 611.850 1321.025 612.130 1325.025 ;
        RECT 1759.660 17.410 1759.800 1328.050 ;
        RECT 1759.660 17.270 1763.020 17.410 ;
        RECT 1762.880 2.400 1763.020 17.270 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 698.350 205.260 698.670 205.320 ;
        RECT 1780.270 205.260 1780.590 205.320 ;
        RECT 698.350 205.120 1780.590 205.260 ;
        RECT 698.350 205.060 698.670 205.120 ;
        RECT 1780.270 205.060 1780.590 205.120 ;
      LAYER via ;
        RECT 698.380 205.060 698.640 205.320 ;
        RECT 1780.300 205.060 1780.560 205.320 ;
      LAYER met2 ;
        RECT 698.330 216.000 698.610 220.000 ;
        RECT 698.440 205.350 698.580 216.000 ;
        RECT 698.380 205.030 698.640 205.350 ;
        RECT 1780.300 205.030 1780.560 205.350 ;
        RECT 1780.360 17.410 1780.500 205.030 ;
        RECT 1780.360 17.270 1780.960 17.410 ;
        RECT 1780.820 2.400 1780.960 17.270 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 372.880 1421.330 372.940 ;
        RECT 1794.070 372.880 1794.390 372.940 ;
        RECT 1421.010 372.740 1794.390 372.880 ;
        RECT 1421.010 372.680 1421.330 372.740 ;
        RECT 1794.070 372.680 1794.390 372.740 ;
      LAYER via ;
        RECT 1421.040 372.680 1421.300 372.940 ;
        RECT 1794.100 372.680 1794.360 372.940 ;
      LAYER met2 ;
        RECT 1421.030 372.795 1421.310 373.165 ;
        RECT 1421.040 372.650 1421.300 372.795 ;
        RECT 1794.100 372.650 1794.360 372.970 ;
        RECT 1794.160 17.410 1794.300 372.650 ;
        RECT 1794.160 17.270 1798.900 17.410 ;
        RECT 1798.760 2.400 1798.900 17.270 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
      LAYER via2 ;
        RECT 1421.030 372.840 1421.310 373.120 ;
      LAYER met3 ;
        RECT 1421.005 373.130 1421.335 373.145 ;
        RECT 1408.060 373.040 1421.335 373.130 ;
        RECT 1404.305 372.830 1421.335 373.040 ;
        RECT 1404.305 372.440 1408.305 372.830 ;
        RECT 1421.005 372.815 1421.335 372.830 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 307.350 217.160 307.670 217.220 ;
        RECT 1814.770 217.160 1815.090 217.220 ;
        RECT 307.350 217.020 1815.090 217.160 ;
        RECT 307.350 216.960 307.670 217.020 ;
        RECT 1814.770 216.960 1815.090 217.020 ;
      LAYER via ;
        RECT 307.380 216.960 307.640 217.220 ;
        RECT 1814.800 216.960 1815.060 217.220 ;
      LAYER met2 ;
        RECT 307.370 292.555 307.650 292.925 ;
        RECT 307.440 217.250 307.580 292.555 ;
        RECT 307.380 216.930 307.640 217.250 ;
        RECT 1814.800 216.930 1815.060 217.250 ;
        RECT 1814.860 17.410 1815.000 216.930 ;
        RECT 1814.860 17.270 1816.840 17.410 ;
        RECT 1816.700 2.400 1816.840 17.270 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
      LAYER via2 ;
        RECT 307.370 292.600 307.650 292.880 ;
      LAYER met3 ;
        RECT 307.345 292.890 307.675 292.905 ;
        RECT 307.345 292.800 310.500 292.890 ;
        RECT 307.345 292.590 314.000 292.800 ;
        RECT 307.345 292.575 307.675 292.590 ;
        RECT 310.000 292.200 314.000 292.590 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1286.230 206.280 1286.550 206.340 ;
        RECT 1828.570 206.280 1828.890 206.340 ;
        RECT 1286.230 206.140 1828.890 206.280 ;
        RECT 1286.230 206.080 1286.550 206.140 ;
        RECT 1828.570 206.080 1828.890 206.140 ;
        RECT 1828.570 16.900 1828.890 16.960 ;
        RECT 1834.550 16.900 1834.870 16.960 ;
        RECT 1828.570 16.760 1834.870 16.900 ;
        RECT 1828.570 16.700 1828.890 16.760 ;
        RECT 1834.550 16.700 1834.870 16.760 ;
      LAYER via ;
        RECT 1286.260 206.080 1286.520 206.340 ;
        RECT 1828.600 206.080 1828.860 206.340 ;
        RECT 1828.600 16.700 1828.860 16.960 ;
        RECT 1834.580 16.700 1834.840 16.960 ;
      LAYER met2 ;
        RECT 1286.210 216.000 1286.490 220.000 ;
        RECT 1286.320 206.370 1286.460 216.000 ;
        RECT 1286.260 206.050 1286.520 206.370 ;
        RECT 1828.600 206.050 1828.860 206.370 ;
        RECT 1828.660 16.990 1828.800 206.050 ;
        RECT 1828.600 16.670 1828.860 16.990 ;
        RECT 1834.580 16.670 1834.840 16.990 ;
        RECT 1834.640 2.400 1834.780 16.670 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 721.810 1321.280 722.130 1321.540 ;
        RECT 721.900 1320.120 722.040 1321.280 ;
        RECT 1849.270 1320.120 1849.590 1320.180 ;
        RECT 721.900 1319.980 1849.590 1320.120 ;
        RECT 1849.270 1319.920 1849.590 1319.980 ;
      LAYER via ;
        RECT 721.840 1321.280 722.100 1321.540 ;
        RECT 1849.300 1319.920 1849.560 1320.180 ;
      LAYER met2 ;
        RECT 720.410 1321.650 720.690 1325.025 ;
        RECT 720.410 1321.570 722.040 1321.650 ;
        RECT 720.410 1321.510 722.100 1321.570 ;
        RECT 720.410 1321.025 720.690 1321.510 ;
        RECT 721.840 1321.250 722.100 1321.510 ;
        RECT 1849.300 1319.890 1849.560 1320.210 ;
        RECT 1849.360 17.410 1849.500 1319.890 ;
        RECT 1849.360 17.270 1852.260 17.410 ;
        RECT 1852.120 2.400 1852.260 17.270 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1420.090 531.660 1420.410 531.720 ;
        RECT 1870.430 531.660 1870.750 531.720 ;
        RECT 1420.090 531.520 1870.750 531.660 ;
        RECT 1420.090 531.460 1420.410 531.520 ;
        RECT 1870.430 531.460 1870.750 531.520 ;
      LAYER via ;
        RECT 1420.120 531.460 1420.380 531.720 ;
        RECT 1870.460 531.460 1870.720 531.720 ;
      LAYER met2 ;
        RECT 1420.110 534.635 1420.390 535.005 ;
        RECT 1420.180 531.750 1420.320 534.635 ;
        RECT 1420.120 531.430 1420.380 531.750 ;
        RECT 1870.460 531.430 1870.720 531.750 ;
        RECT 1870.520 7.210 1870.660 531.430 ;
        RECT 1870.060 7.070 1870.660 7.210 ;
        RECT 1870.060 2.400 1870.200 7.070 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
      LAYER via2 ;
        RECT 1420.110 534.680 1420.390 534.960 ;
      LAYER met3 ;
        RECT 1420.085 534.970 1420.415 534.985 ;
        RECT 1408.060 534.880 1420.415 534.970 ;
        RECT 1404.305 534.670 1420.415 534.880 ;
        RECT 1404.305 534.280 1408.305 534.670 ;
        RECT 1420.085 534.655 1420.415 534.670 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 745.345 186.405 745.515 218.875 ;
        RECT 745.345 89.845 745.515 137.955 ;
      LAYER mcon ;
        RECT 745.345 218.705 745.515 218.875 ;
        RECT 745.345 137.785 745.515 137.955 ;
      LAYER met1 ;
        RECT 305.050 218.860 305.370 218.920 ;
        RECT 745.285 218.860 745.575 218.905 ;
        RECT 305.050 218.720 745.575 218.860 ;
        RECT 305.050 218.660 305.370 218.720 ;
        RECT 745.285 218.675 745.575 218.720 ;
        RECT 745.270 186.560 745.590 186.620 ;
        RECT 745.075 186.420 745.590 186.560 ;
        RECT 745.270 186.360 745.590 186.420 ;
        RECT 745.270 137.940 745.590 138.000 ;
        RECT 745.075 137.800 745.590 137.940 ;
        RECT 745.270 137.740 745.590 137.800 ;
        RECT 745.270 90.000 745.590 90.060 ;
        RECT 745.075 89.860 745.590 90.000 ;
        RECT 745.270 89.800 745.590 89.860 ;
        RECT 745.270 62.260 745.590 62.520 ;
        RECT 745.360 61.440 745.500 62.260 ;
        RECT 746.190 61.440 746.510 61.500 ;
        RECT 745.360 61.300 746.510 61.440 ;
        RECT 746.190 61.240 746.510 61.300 ;
      LAYER via ;
        RECT 305.080 218.660 305.340 218.920 ;
        RECT 745.300 186.360 745.560 186.620 ;
        RECT 745.300 137.740 745.560 138.000 ;
        RECT 745.300 89.800 745.560 90.060 ;
        RECT 745.300 62.260 745.560 62.520 ;
        RECT 746.220 61.240 746.480 61.500 ;
      LAYER met2 ;
        RECT 305.070 351.035 305.350 351.405 ;
        RECT 305.140 218.950 305.280 351.035 ;
        RECT 305.080 218.630 305.340 218.950 ;
        RECT 745.300 186.330 745.560 186.650 ;
        RECT 745.360 138.030 745.500 186.330 ;
        RECT 745.300 137.710 745.560 138.030 ;
        RECT 745.300 89.770 745.560 90.090 ;
        RECT 745.360 62.550 745.500 89.770 ;
        RECT 745.300 62.230 745.560 62.550 ;
        RECT 746.220 61.210 746.480 61.530 ;
        RECT 746.280 2.400 746.420 61.210 ;
        RECT 746.070 -4.800 746.630 2.400 ;
      LAYER via2 ;
        RECT 305.070 351.080 305.350 351.360 ;
      LAYER met3 ;
        RECT 305.045 351.370 305.375 351.385 ;
        RECT 305.045 351.280 310.500 351.370 ;
        RECT 305.045 351.070 314.000 351.280 ;
        RECT 305.045 351.055 305.375 351.070 ;
        RECT 310.000 350.680 314.000 351.070 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.430 203.560 559.750 203.620 ;
        RECT 1883.770 203.560 1884.090 203.620 ;
        RECT 559.430 203.420 1884.090 203.560 ;
        RECT 559.430 203.360 559.750 203.420 ;
        RECT 1883.770 203.360 1884.090 203.420 ;
      LAYER via ;
        RECT 559.460 203.360 559.720 203.620 ;
        RECT 1883.800 203.360 1884.060 203.620 ;
      LAYER met2 ;
        RECT 559.410 216.000 559.690 220.000 ;
        RECT 559.520 203.650 559.660 216.000 ;
        RECT 559.460 203.330 559.720 203.650 ;
        RECT 1883.800 203.330 1884.060 203.650 ;
        RECT 1883.860 17.410 1884.000 203.330 ;
        RECT 1883.860 17.270 1888.140 17.410 ;
        RECT 1888.000 2.400 1888.140 17.270 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1197.910 205.940 1198.230 206.000 ;
        RECT 1904.470 205.940 1904.790 206.000 ;
        RECT 1197.910 205.800 1904.790 205.940 ;
        RECT 1197.910 205.740 1198.230 205.800 ;
        RECT 1904.470 205.740 1904.790 205.800 ;
      LAYER via ;
        RECT 1197.940 205.740 1198.200 206.000 ;
        RECT 1904.500 205.740 1904.760 206.000 ;
      LAYER met2 ;
        RECT 1197.890 216.000 1198.170 220.000 ;
        RECT 1198.000 206.030 1198.140 216.000 ;
        RECT 1197.940 205.710 1198.200 206.030 ;
        RECT 1904.500 205.710 1904.760 206.030 ;
        RECT 1904.560 17.410 1904.700 205.710 ;
        RECT 1904.560 17.270 1906.080 17.410 ;
        RECT 1905.940 2.400 1906.080 17.270 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 767.350 204.920 767.670 204.980 ;
        RECT 1918.270 204.920 1918.590 204.980 ;
        RECT 767.350 204.780 1918.590 204.920 ;
        RECT 767.350 204.720 767.670 204.780 ;
        RECT 1918.270 204.720 1918.590 204.780 ;
      LAYER via ;
        RECT 767.380 204.720 767.640 204.980 ;
        RECT 1918.300 204.720 1918.560 204.980 ;
      LAYER met2 ;
        RECT 767.330 216.000 767.610 220.000 ;
        RECT 767.440 205.010 767.580 216.000 ;
        RECT 767.380 204.690 767.640 205.010 ;
        RECT 1918.300 204.690 1918.560 205.010 ;
        RECT 1918.360 17.410 1918.500 204.690 ;
        RECT 1918.360 17.270 1923.560 17.410 ;
        RECT 1923.420 2.400 1923.560 17.270 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1255.410 33.560 1255.730 33.620 ;
        RECT 1941.270 33.560 1941.590 33.620 ;
        RECT 1255.410 33.420 1941.590 33.560 ;
        RECT 1255.410 33.360 1255.730 33.420 ;
        RECT 1941.270 33.360 1941.590 33.420 ;
      LAYER via ;
        RECT 1255.440 33.360 1255.700 33.620 ;
        RECT 1941.300 33.360 1941.560 33.620 ;
      LAYER met2 ;
        RECT 1252.170 216.650 1252.450 220.000 ;
        RECT 1252.170 216.510 1255.640 216.650 ;
        RECT 1252.170 216.000 1252.450 216.510 ;
        RECT 1255.500 33.650 1255.640 216.510 ;
        RECT 1255.440 33.330 1255.700 33.650 ;
        RECT 1941.300 33.330 1941.560 33.650 ;
        RECT 1941.360 2.400 1941.500 33.330 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 298.610 196.760 298.930 196.820 ;
        RECT 1953.230 196.760 1953.550 196.820 ;
        RECT 298.610 196.620 1953.550 196.760 ;
        RECT 298.610 196.560 298.930 196.620 ;
        RECT 1953.230 196.560 1953.550 196.620 ;
        RECT 1953.230 19.620 1953.550 19.680 ;
        RECT 1959.210 19.620 1959.530 19.680 ;
        RECT 1953.230 19.480 1959.530 19.620 ;
        RECT 1953.230 19.420 1953.550 19.480 ;
        RECT 1959.210 19.420 1959.530 19.480 ;
      LAYER via ;
        RECT 298.640 196.560 298.900 196.820 ;
        RECT 1953.260 196.560 1953.520 196.820 ;
        RECT 1953.260 19.420 1953.520 19.680 ;
        RECT 1959.240 19.420 1959.500 19.680 ;
      LAYER met2 ;
        RECT 298.630 439.435 298.910 439.805 ;
        RECT 298.700 196.850 298.840 439.435 ;
        RECT 298.640 196.530 298.900 196.850 ;
        RECT 1953.260 196.530 1953.520 196.850 ;
        RECT 1953.320 19.710 1953.460 196.530 ;
        RECT 1953.260 19.390 1953.520 19.710 ;
        RECT 1959.240 19.390 1959.500 19.710 ;
        RECT 1959.300 2.400 1959.440 19.390 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
      LAYER via2 ;
        RECT 298.630 439.480 298.910 439.760 ;
      LAYER met3 ;
        RECT 298.605 439.770 298.935 439.785 ;
        RECT 298.605 439.680 310.500 439.770 ;
        RECT 298.605 439.470 314.000 439.680 ;
        RECT 298.605 439.455 298.935 439.470 ;
        RECT 310.000 439.080 314.000 439.470 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 924.210 39.340 924.530 39.400 ;
        RECT 1977.150 39.340 1977.470 39.400 ;
        RECT 924.210 39.200 1977.470 39.340 ;
        RECT 924.210 39.140 924.530 39.200 ;
        RECT 1977.150 39.140 1977.470 39.200 ;
      LAYER via ;
        RECT 924.240 39.140 924.500 39.400 ;
        RECT 1977.180 39.140 1977.440 39.400 ;
      LAYER met2 ;
        RECT 920.970 216.650 921.250 220.000 ;
        RECT 920.970 216.510 924.440 216.650 ;
        RECT 920.970 216.000 921.250 216.510 ;
        RECT 924.300 39.430 924.440 216.510 ;
        RECT 924.240 39.110 924.500 39.430 ;
        RECT 1977.180 39.110 1977.440 39.430 ;
        RECT 1977.240 2.400 1977.380 39.110 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 317.470 200.500 317.790 200.560 ;
        RECT 327.590 200.500 327.910 200.560 ;
        RECT 317.470 200.360 327.910 200.500 ;
        RECT 317.470 200.300 317.790 200.360 ;
        RECT 327.590 200.300 327.910 200.360 ;
        RECT 327.590 38.320 327.910 38.380 ;
        RECT 1995.090 38.320 1995.410 38.380 ;
        RECT 327.590 38.180 1995.410 38.320 ;
        RECT 327.590 38.120 327.910 38.180 ;
        RECT 1995.090 38.120 1995.410 38.180 ;
      LAYER via ;
        RECT 317.500 200.300 317.760 200.560 ;
        RECT 327.620 200.300 327.880 200.560 ;
        RECT 327.620 38.120 327.880 38.380 ;
        RECT 1995.120 38.120 1995.380 38.380 ;
      LAYER met2 ;
        RECT 317.450 216.000 317.730 220.000 ;
        RECT 317.560 200.590 317.700 216.000 ;
        RECT 317.500 200.270 317.760 200.590 ;
        RECT 327.620 200.270 327.880 200.590 ;
        RECT 327.680 38.410 327.820 200.270 ;
        RECT 327.620 38.090 327.880 38.410 ;
        RECT 1995.120 38.090 1995.380 38.410 ;
        RECT 1995.180 2.400 1995.320 38.090 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1076.010 121.280 1076.330 121.340 ;
        RECT 2007.970 121.280 2008.290 121.340 ;
        RECT 1076.010 121.140 2008.290 121.280 ;
        RECT 1076.010 121.080 1076.330 121.140 ;
        RECT 2007.970 121.080 2008.290 121.140 ;
        RECT 2007.970 2.960 2008.290 3.020 ;
        RECT 2012.570 2.960 2012.890 3.020 ;
        RECT 2007.970 2.820 2012.890 2.960 ;
        RECT 2007.970 2.760 2008.290 2.820 ;
        RECT 2012.570 2.760 2012.890 2.820 ;
      LAYER via ;
        RECT 1076.040 121.080 1076.300 121.340 ;
        RECT 2008.000 121.080 2008.260 121.340 ;
        RECT 2008.000 2.760 2008.260 3.020 ;
        RECT 2012.600 2.760 2012.860 3.020 ;
      LAYER met2 ;
        RECT 1073.690 216.650 1073.970 220.000 ;
        RECT 1073.690 216.510 1076.240 216.650 ;
        RECT 1073.690 216.000 1073.970 216.510 ;
        RECT 1076.100 121.370 1076.240 216.510 ;
        RECT 1076.040 121.050 1076.300 121.370 ;
        RECT 2008.000 121.050 2008.260 121.370 ;
        RECT 2008.060 3.050 2008.200 121.050 ;
        RECT 2008.000 2.730 2008.260 3.050 ;
        RECT 2012.600 2.730 2012.860 3.050 ;
        RECT 2012.660 2.400 2012.800 2.730 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1173.070 205.600 1173.390 205.660 ;
        RECT 2028.670 205.600 2028.990 205.660 ;
        RECT 1173.070 205.460 2028.990 205.600 ;
        RECT 1173.070 205.400 1173.390 205.460 ;
        RECT 2028.670 205.400 2028.990 205.460 ;
      LAYER via ;
        RECT 1173.100 205.400 1173.360 205.660 ;
        RECT 2028.700 205.400 2028.960 205.660 ;
      LAYER met2 ;
        RECT 1173.050 216.000 1173.330 220.000 ;
        RECT 1173.160 205.690 1173.300 216.000 ;
        RECT 1173.100 205.370 1173.360 205.690 ;
        RECT 2028.700 205.370 2028.960 205.690 ;
        RECT 2028.760 16.730 2028.900 205.370 ;
        RECT 2028.760 16.590 2030.740 16.730 ;
        RECT 2030.600 2.400 2030.740 16.590 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1066.350 1341.540 1066.670 1341.600 ;
        RECT 2042.470 1341.540 2042.790 1341.600 ;
        RECT 1066.350 1341.400 2042.790 1341.540 ;
        RECT 1066.350 1341.340 1066.670 1341.400 ;
        RECT 2042.470 1341.340 2042.790 1341.400 ;
        RECT 2042.470 19.620 2042.790 19.680 ;
        RECT 2048.450 19.620 2048.770 19.680 ;
        RECT 2042.470 19.480 2048.770 19.620 ;
        RECT 2042.470 19.420 2042.790 19.480 ;
        RECT 2048.450 19.420 2048.770 19.480 ;
      LAYER via ;
        RECT 1066.380 1341.340 1066.640 1341.600 ;
        RECT 2042.500 1341.340 2042.760 1341.600 ;
        RECT 2042.500 19.420 2042.760 19.680 ;
        RECT 2048.480 19.420 2048.740 19.680 ;
      LAYER met2 ;
        RECT 1066.380 1341.310 1066.640 1341.630 ;
        RECT 2042.500 1341.310 2042.760 1341.630 ;
        RECT 1066.440 1325.025 1066.580 1341.310 ;
        RECT 1066.330 1321.025 1066.610 1325.025 ;
        RECT 2042.560 19.710 2042.700 1341.310 ;
        RECT 2042.500 19.390 2042.760 19.710 ;
        RECT 2048.480 19.390 2048.740 19.710 ;
        RECT 2048.540 2.400 2048.680 19.390 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 763.745 2.805 763.915 14.195 ;
      LAYER mcon ;
        RECT 763.745 14.025 763.915 14.195 ;
      LAYER met1 ;
        RECT 763.685 14.180 763.975 14.225 ;
        RECT 765.510 14.180 765.830 14.240 ;
        RECT 763.685 14.040 765.830 14.180 ;
        RECT 763.685 13.995 763.975 14.040 ;
        RECT 765.510 13.980 765.830 14.040 ;
        RECT 763.670 2.960 763.990 3.020 ;
        RECT 763.475 2.820 763.990 2.960 ;
        RECT 763.670 2.760 763.990 2.820 ;
      LAYER via ;
        RECT 765.540 13.980 765.800 14.240 ;
        RECT 763.700 2.760 763.960 3.020 ;
      LAYER met2 ;
        RECT 997.370 1346.555 997.650 1346.925 ;
        RECT 997.440 1325.025 997.580 1346.555 ;
        RECT 997.330 1321.025 997.610 1325.025 ;
        RECT 765.530 210.955 765.810 211.325 ;
        RECT 765.600 14.270 765.740 210.955 ;
        RECT 765.540 13.950 765.800 14.270 ;
        RECT 763.700 2.730 763.960 3.050 ;
        RECT 763.760 2.400 763.900 2.730 ;
        RECT 763.550 -4.800 764.110 2.400 ;
      LAYER via2 ;
        RECT 997.370 1346.600 997.650 1346.880 ;
        RECT 765.530 211.000 765.810 211.280 ;
      LAYER met3 ;
        RECT 997.345 1346.890 997.675 1346.905 ;
        RECT 1412.470 1346.890 1412.850 1346.900 ;
        RECT 997.345 1346.590 1412.850 1346.890 ;
        RECT 997.345 1346.575 997.675 1346.590 ;
        RECT 1412.470 1346.580 1412.850 1346.590 ;
        RECT 765.505 211.290 765.835 211.305 ;
        RECT 1384.870 211.290 1385.250 211.300 ;
        RECT 765.505 210.990 1385.250 211.290 ;
        RECT 765.505 210.975 765.835 210.990 ;
        RECT 1384.870 210.980 1385.250 210.990 ;
      LAYER via3 ;
        RECT 1412.500 1346.580 1412.820 1346.900 ;
        RECT 1384.900 210.980 1385.220 211.300 ;
      LAYER met4 ;
        RECT 1412.495 1346.575 1412.825 1346.905 ;
        RECT 1412.510 223.290 1412.810 1346.575 ;
        RECT 1384.470 222.110 1385.650 223.290 ;
        RECT 1412.070 222.110 1413.250 223.290 ;
        RECT 1384.910 211.305 1385.210 222.110 ;
        RECT 1384.895 210.975 1385.225 211.305 ;
      LAYER met5 ;
        RECT 1384.260 221.900 1413.460 223.500 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 908.110 1347.660 908.430 1347.720 ;
        RECT 2063.170 1347.660 2063.490 1347.720 ;
        RECT 908.110 1347.520 2063.490 1347.660 ;
        RECT 908.110 1347.460 908.430 1347.520 ;
        RECT 2063.170 1347.460 2063.490 1347.520 ;
        RECT 2063.170 2.960 2063.490 3.020 ;
        RECT 2066.390 2.960 2066.710 3.020 ;
        RECT 2063.170 2.820 2066.710 2.960 ;
        RECT 2063.170 2.760 2063.490 2.820 ;
        RECT 2066.390 2.760 2066.710 2.820 ;
      LAYER via ;
        RECT 908.140 1347.460 908.400 1347.720 ;
        RECT 2063.200 1347.460 2063.460 1347.720 ;
        RECT 2063.200 2.760 2063.460 3.020 ;
        RECT 2066.420 2.760 2066.680 3.020 ;
      LAYER met2 ;
        RECT 908.140 1347.430 908.400 1347.750 ;
        RECT 2063.200 1347.430 2063.460 1347.750 ;
        RECT 908.200 1325.025 908.340 1347.430 ;
        RECT 908.090 1321.025 908.370 1325.025 ;
        RECT 2063.260 3.050 2063.400 1347.430 ;
        RECT 2063.200 2.730 2063.460 3.050 ;
        RECT 2066.420 2.730 2066.680 3.050 ;
        RECT 2066.480 2.400 2066.620 2.730 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 695.590 1346.980 695.910 1347.040 ;
        RECT 2084.330 1346.980 2084.650 1347.040 ;
        RECT 695.590 1346.840 2084.650 1346.980 ;
        RECT 695.590 1346.780 695.910 1346.840 ;
        RECT 2084.330 1346.780 2084.650 1346.840 ;
      LAYER via ;
        RECT 695.620 1346.780 695.880 1347.040 ;
        RECT 2084.360 1346.780 2084.620 1347.040 ;
      LAYER met2 ;
        RECT 695.620 1346.750 695.880 1347.070 ;
        RECT 2084.360 1346.750 2084.620 1347.070 ;
        RECT 695.680 1325.025 695.820 1346.750 ;
        RECT 695.570 1321.025 695.850 1325.025 ;
        RECT 2084.420 2.400 2084.560 1346.750 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 562.190 1346.300 562.510 1346.360 ;
        RECT 2097.670 1346.300 2097.990 1346.360 ;
        RECT 562.190 1346.160 2097.990 1346.300 ;
        RECT 562.190 1346.100 562.510 1346.160 ;
        RECT 2097.670 1346.100 2097.990 1346.160 ;
        RECT 2097.670 2.960 2097.990 3.020 ;
        RECT 2101.810 2.960 2102.130 3.020 ;
        RECT 2097.670 2.820 2102.130 2.960 ;
        RECT 2097.670 2.760 2097.990 2.820 ;
        RECT 2101.810 2.760 2102.130 2.820 ;
      LAYER via ;
        RECT 562.220 1346.100 562.480 1346.360 ;
        RECT 2097.700 1346.100 2097.960 1346.360 ;
        RECT 2097.700 2.760 2097.960 3.020 ;
        RECT 2101.840 2.760 2102.100 3.020 ;
      LAYER met2 ;
        RECT 562.220 1346.070 562.480 1346.390 ;
        RECT 2097.700 1346.070 2097.960 1346.390 ;
        RECT 562.280 1325.025 562.420 1346.070 ;
        RECT 562.170 1321.025 562.450 1325.025 ;
        RECT 2097.760 3.050 2097.900 1346.070 ;
        RECT 2097.700 2.730 2097.960 3.050 ;
        RECT 2101.840 2.730 2102.100 3.050 ;
        RECT 2101.900 2.400 2102.040 2.730 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1420.090 545.260 1420.410 545.320 ;
        RECT 2118.370 545.260 2118.690 545.320 ;
        RECT 1420.090 545.120 2118.690 545.260 ;
        RECT 1420.090 545.060 1420.410 545.120 ;
        RECT 2118.370 545.060 2118.690 545.120 ;
      LAYER via ;
        RECT 1420.120 545.060 1420.380 545.320 ;
        RECT 2118.400 545.060 2118.660 545.320 ;
      LAYER met2 ;
        RECT 1420.110 548.235 1420.390 548.605 ;
        RECT 1420.180 545.350 1420.320 548.235 ;
        RECT 1420.120 545.030 1420.380 545.350 ;
        RECT 2118.400 545.030 2118.660 545.350 ;
        RECT 2118.460 17.410 2118.600 545.030 ;
        RECT 2118.460 17.270 2119.980 17.410 ;
        RECT 2119.840 2.400 2119.980 17.270 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
      LAYER via2 ;
        RECT 1420.110 548.280 1420.390 548.560 ;
      LAYER met3 ;
        RECT 1420.085 548.570 1420.415 548.585 ;
        RECT 1408.060 548.480 1420.415 548.570 ;
        RECT 1404.305 548.270 1420.415 548.480 ;
        RECT 1404.305 547.880 1408.305 548.270 ;
        RECT 1420.085 548.255 1420.415 548.270 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1418.710 683.300 1419.030 683.360 ;
        RECT 2132.170 683.300 2132.490 683.360 ;
        RECT 1418.710 683.160 2132.490 683.300 ;
        RECT 1418.710 683.100 1419.030 683.160 ;
        RECT 2132.170 683.100 2132.490 683.160 ;
      LAYER via ;
        RECT 1418.740 683.100 1419.000 683.360 ;
        RECT 2132.200 683.100 2132.460 683.360 ;
      LAYER met2 ;
        RECT 1418.730 688.315 1419.010 688.685 ;
        RECT 1418.800 683.390 1418.940 688.315 ;
        RECT 1418.740 683.070 1419.000 683.390 ;
        RECT 2132.200 683.070 2132.460 683.390 ;
        RECT 2132.260 17.410 2132.400 683.070 ;
        RECT 2132.260 17.270 2137.920 17.410 ;
        RECT 2137.780 2.400 2137.920 17.270 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
      LAYER via2 ;
        RECT 1418.730 688.360 1419.010 688.640 ;
      LAYER met3 ;
        RECT 1418.705 688.650 1419.035 688.665 ;
        RECT 1408.060 688.560 1419.035 688.650 ;
        RECT 1404.305 688.350 1419.035 688.560 ;
        RECT 1404.305 687.960 1408.305 688.350 ;
        RECT 1418.705 688.335 1419.035 688.350 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 993.720 1421.330 993.780 ;
        RECT 2152.870 993.720 2153.190 993.780 ;
        RECT 1421.010 993.580 2153.190 993.720 ;
        RECT 1421.010 993.520 1421.330 993.580 ;
        RECT 2152.870 993.520 2153.190 993.580 ;
      LAYER via ;
        RECT 1421.040 993.520 1421.300 993.780 ;
        RECT 2152.900 993.520 2153.160 993.780 ;
      LAYER met2 ;
        RECT 1421.030 994.315 1421.310 994.685 ;
        RECT 1421.100 993.810 1421.240 994.315 ;
        RECT 1421.040 993.490 1421.300 993.810 ;
        RECT 2152.900 993.490 2153.160 993.810 ;
        RECT 2152.960 17.410 2153.100 993.490 ;
        RECT 2152.960 17.270 2155.860 17.410 ;
        RECT 2155.720 2.400 2155.860 17.270 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
      LAYER via2 ;
        RECT 1421.030 994.360 1421.310 994.640 ;
      LAYER met3 ;
        RECT 1421.005 994.650 1421.335 994.665 ;
        RECT 1408.060 994.560 1421.335 994.650 ;
        RECT 1404.305 994.350 1421.335 994.560 ;
        RECT 1404.305 993.960 1408.305 994.350 ;
        RECT 1421.005 994.335 1421.335 994.350 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1418.710 559.200 1419.030 559.260 ;
        RECT 2166.670 559.200 2166.990 559.260 ;
        RECT 1418.710 559.060 2166.990 559.200 ;
        RECT 1418.710 559.000 1419.030 559.060 ;
        RECT 2166.670 559.000 2166.990 559.060 ;
        RECT 2166.670 17.580 2166.990 17.640 ;
        RECT 2173.110 17.580 2173.430 17.640 ;
        RECT 2166.670 17.440 2173.430 17.580 ;
        RECT 2166.670 17.380 2166.990 17.440 ;
        RECT 2173.110 17.380 2173.430 17.440 ;
      LAYER via ;
        RECT 1418.740 559.000 1419.000 559.260 ;
        RECT 2166.700 559.000 2166.960 559.260 ;
        RECT 2166.700 17.380 2166.960 17.640 ;
        RECT 2173.140 17.380 2173.400 17.640 ;
      LAYER met2 ;
        RECT 1418.730 563.195 1419.010 563.565 ;
        RECT 1418.800 559.290 1418.940 563.195 ;
        RECT 1418.740 558.970 1419.000 559.290 ;
        RECT 2166.700 558.970 2166.960 559.290 ;
        RECT 2166.760 17.670 2166.900 558.970 ;
        RECT 2166.700 17.350 2166.960 17.670 ;
        RECT 2173.140 17.350 2173.400 17.670 ;
        RECT 2173.200 2.400 2173.340 17.350 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
      LAYER via2 ;
        RECT 1418.730 563.240 1419.010 563.520 ;
      LAYER met3 ;
        RECT 1418.705 563.530 1419.035 563.545 ;
        RECT 1408.060 563.440 1419.035 563.530 ;
        RECT 1404.305 563.230 1419.035 563.440 ;
        RECT 1404.305 562.840 1408.305 563.230 ;
        RECT 1418.705 563.215 1419.035 563.230 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 859.350 1326.240 859.670 1326.300 ;
        RECT 2187.370 1326.240 2187.690 1326.300 ;
        RECT 859.350 1326.100 2187.690 1326.240 ;
        RECT 859.350 1326.040 859.670 1326.100 ;
        RECT 2187.370 1326.040 2187.690 1326.100 ;
      LAYER via ;
        RECT 859.380 1326.040 859.640 1326.300 ;
        RECT 2187.400 1326.040 2187.660 1326.300 ;
      LAYER met2 ;
        RECT 859.380 1326.010 859.640 1326.330 ;
        RECT 2187.400 1326.010 2187.660 1326.330 ;
        RECT 859.440 1325.025 859.580 1326.010 ;
        RECT 859.330 1321.025 859.610 1325.025 ;
        RECT 2187.460 17.410 2187.600 1326.010 ;
        RECT 2187.460 17.270 2191.280 17.410 ;
        RECT 2191.140 2.400 2191.280 17.270 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1227.350 204.580 1227.670 204.640 ;
        RECT 2208.070 204.580 2208.390 204.640 ;
        RECT 1227.350 204.440 2208.390 204.580 ;
        RECT 1227.350 204.380 1227.670 204.440 ;
        RECT 2208.070 204.380 2208.390 204.440 ;
      LAYER via ;
        RECT 1227.380 204.380 1227.640 204.640 ;
        RECT 2208.100 204.380 2208.360 204.640 ;
      LAYER met2 ;
        RECT 1227.330 216.000 1227.610 220.000 ;
        RECT 1227.440 204.670 1227.580 216.000 ;
        RECT 1227.380 204.350 1227.640 204.670 ;
        RECT 2208.100 204.350 2208.360 204.670 ;
        RECT 2208.160 17.410 2208.300 204.350 ;
        RECT 2208.160 17.270 2209.220 17.410 ;
        RECT 2209.080 2.400 2209.220 17.270 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 293.090 58.720 293.410 58.780 ;
        RECT 2221.870 58.720 2222.190 58.780 ;
        RECT 293.090 58.580 2222.190 58.720 ;
        RECT 293.090 58.520 293.410 58.580 ;
        RECT 2221.870 58.520 2222.190 58.580 ;
      LAYER via ;
        RECT 293.120 58.520 293.380 58.780 ;
        RECT 2221.900 58.520 2222.160 58.780 ;
      LAYER met2 ;
        RECT 293.110 599.915 293.390 600.285 ;
        RECT 293.180 58.810 293.320 599.915 ;
        RECT 293.120 58.490 293.380 58.810 ;
        RECT 2221.900 58.490 2222.160 58.810 ;
        RECT 2221.960 17.410 2222.100 58.490 ;
        RECT 2221.960 17.270 2227.160 17.410 ;
        RECT 2227.020 2.400 2227.160 17.270 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
      LAYER via2 ;
        RECT 293.110 599.960 293.390 600.240 ;
      LAYER met3 ;
        RECT 293.085 600.250 293.415 600.265 ;
        RECT 293.085 600.160 310.500 600.250 ;
        RECT 293.085 599.950 314.000 600.160 ;
        RECT 293.085 599.935 293.415 599.950 ;
        RECT 310.000 599.560 314.000 599.950 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 503.780 1421.330 503.840 ;
        RECT 1431.130 503.780 1431.450 503.840 ;
        RECT 1421.010 503.640 1431.450 503.780 ;
        RECT 1421.010 503.580 1421.330 503.640 ;
        RECT 1431.130 503.580 1431.450 503.640 ;
        RECT 786.210 211.720 786.530 211.780 ;
        RECT 1431.130 211.720 1431.450 211.780 ;
        RECT 786.210 211.580 1431.450 211.720 ;
        RECT 786.210 211.520 786.530 211.580 ;
        RECT 1431.130 211.520 1431.450 211.580 ;
        RECT 781.610 16.900 781.930 16.960 ;
        RECT 786.210 16.900 786.530 16.960 ;
        RECT 781.610 16.760 786.530 16.900 ;
        RECT 781.610 16.700 781.930 16.760 ;
        RECT 786.210 16.700 786.530 16.760 ;
      LAYER via ;
        RECT 1421.040 503.580 1421.300 503.840 ;
        RECT 1431.160 503.580 1431.420 503.840 ;
        RECT 786.240 211.520 786.500 211.780 ;
        RECT 1431.160 211.520 1431.420 211.780 ;
        RECT 781.640 16.700 781.900 16.960 ;
        RECT 786.240 16.700 786.500 16.960 ;
      LAYER met2 ;
        RECT 1421.030 504.715 1421.310 505.085 ;
        RECT 1421.100 503.870 1421.240 504.715 ;
        RECT 1421.040 503.550 1421.300 503.870 ;
        RECT 1431.160 503.550 1431.420 503.870 ;
        RECT 1431.220 211.810 1431.360 503.550 ;
        RECT 786.240 211.490 786.500 211.810 ;
        RECT 1431.160 211.490 1431.420 211.810 ;
        RECT 786.300 16.990 786.440 211.490 ;
        RECT 781.640 16.670 781.900 16.990 ;
        RECT 786.240 16.670 786.500 16.990 ;
        RECT 781.700 2.400 781.840 16.670 ;
        RECT 781.490 -4.800 782.050 2.400 ;
      LAYER via2 ;
        RECT 1421.030 504.760 1421.310 505.040 ;
      LAYER met3 ;
        RECT 1421.005 505.050 1421.335 505.065 ;
        RECT 1408.060 504.960 1421.335 505.050 ;
        RECT 1404.305 504.750 1421.335 504.960 ;
        RECT 1404.305 504.360 1408.305 504.750 ;
        RECT 1421.005 504.735 1421.335 504.750 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 299.530 169.220 299.850 169.280 ;
        RECT 2242.570 169.220 2242.890 169.280 ;
        RECT 299.530 169.080 2242.890 169.220 ;
        RECT 299.530 169.020 299.850 169.080 ;
        RECT 2242.570 169.020 2242.890 169.080 ;
      LAYER via ;
        RECT 299.560 169.020 299.820 169.280 ;
        RECT 2242.600 169.020 2242.860 169.280 ;
      LAYER met2 ;
        RECT 299.550 322.475 299.830 322.845 ;
        RECT 299.620 169.310 299.760 322.475 ;
        RECT 299.560 168.990 299.820 169.310 ;
        RECT 2242.600 168.990 2242.860 169.310 ;
        RECT 2242.660 17.410 2242.800 168.990 ;
        RECT 2242.660 17.270 2245.100 17.410 ;
        RECT 2244.960 2.400 2245.100 17.270 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
      LAYER via2 ;
        RECT 299.550 322.520 299.830 322.800 ;
      LAYER met3 ;
        RECT 299.525 322.810 299.855 322.825 ;
        RECT 299.525 322.720 310.500 322.810 ;
        RECT 299.525 322.510 314.000 322.720 ;
        RECT 299.525 322.495 299.855 322.510 ;
        RECT 310.000 322.120 314.000 322.510 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1328.550 1335.080 1328.870 1335.140 ;
        RECT 1405.830 1335.080 1406.150 1335.140 ;
        RECT 1328.550 1334.940 1406.150 1335.080 ;
        RECT 1328.550 1334.880 1328.870 1334.940 ;
        RECT 1405.830 1334.880 1406.150 1334.940 ;
        RECT 1405.830 1307.880 1406.150 1307.940 ;
        RECT 2256.830 1307.880 2257.150 1307.940 ;
        RECT 1405.830 1307.740 2257.150 1307.880 ;
        RECT 1405.830 1307.680 1406.150 1307.740 ;
        RECT 2256.830 1307.680 2257.150 1307.740 ;
      LAYER via ;
        RECT 1328.580 1334.880 1328.840 1335.140 ;
        RECT 1405.860 1334.880 1406.120 1335.140 ;
        RECT 1405.860 1307.680 1406.120 1307.940 ;
        RECT 2256.860 1307.680 2257.120 1307.940 ;
      LAYER met2 ;
        RECT 1328.580 1334.850 1328.840 1335.170 ;
        RECT 1405.860 1334.850 1406.120 1335.170 ;
        RECT 1328.640 1325.025 1328.780 1334.850 ;
        RECT 1328.530 1321.025 1328.810 1325.025 ;
        RECT 1405.920 1307.970 1406.060 1334.850 ;
        RECT 1405.860 1307.650 1406.120 1307.970 ;
        RECT 2256.860 1307.650 2257.120 1307.970 ;
        RECT 2256.920 17.410 2257.060 1307.650 ;
        RECT 2256.920 17.270 2262.580 17.410 ;
        RECT 2262.440 2.400 2262.580 17.270 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1388.350 1332.020 1388.670 1332.080 ;
        RECT 1404.450 1332.020 1404.770 1332.080 ;
        RECT 1388.350 1331.880 1404.770 1332.020 ;
        RECT 1388.350 1331.820 1388.670 1331.880 ;
        RECT 1404.450 1331.820 1404.770 1331.880 ;
        RECT 1404.450 1301.080 1404.770 1301.140 ;
        RECT 2277.070 1301.080 2277.390 1301.140 ;
        RECT 1404.450 1300.940 2277.390 1301.080 ;
        RECT 1404.450 1300.880 1404.770 1300.940 ;
        RECT 2277.070 1300.880 2277.390 1300.940 ;
      LAYER via ;
        RECT 1388.380 1331.820 1388.640 1332.080 ;
        RECT 1404.480 1331.820 1404.740 1332.080 ;
        RECT 1404.480 1300.880 1404.740 1301.140 ;
        RECT 2277.100 1300.880 2277.360 1301.140 ;
      LAYER met2 ;
        RECT 1388.380 1331.790 1388.640 1332.110 ;
        RECT 1404.480 1331.790 1404.740 1332.110 ;
        RECT 1388.440 1325.025 1388.580 1331.790 ;
        RECT 1388.330 1321.025 1388.610 1325.025 ;
        RECT 1404.540 1301.170 1404.680 1331.790 ;
        RECT 1404.480 1300.850 1404.740 1301.170 ;
        RECT 2277.100 1300.850 2277.360 1301.170 ;
        RECT 2277.160 17.410 2277.300 1300.850 ;
        RECT 2277.160 17.270 2280.520 17.410 ;
        RECT 2280.380 2.400 2280.520 17.270 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1404.910 1307.540 1405.230 1307.600 ;
        RECT 2297.770 1307.540 2298.090 1307.600 ;
        RECT 1404.910 1307.400 2298.090 1307.540 ;
        RECT 1404.910 1307.340 1405.230 1307.400 ;
        RECT 2297.770 1307.340 2298.090 1307.400 ;
      LAYER via ;
        RECT 1404.940 1307.340 1405.200 1307.600 ;
        RECT 2297.800 1307.340 2298.060 1307.600 ;
      LAYER met2 ;
        RECT 1190.570 1334.995 1190.850 1335.365 ;
        RECT 1405.390 1334.995 1405.670 1335.365 ;
        RECT 1190.640 1325.025 1190.780 1334.995 ;
        RECT 1190.530 1321.025 1190.810 1325.025 ;
        RECT 1405.460 1315.530 1405.600 1334.995 ;
        RECT 1405.000 1315.390 1405.600 1315.530 ;
        RECT 1405.000 1307.630 1405.140 1315.390 ;
        RECT 1404.940 1307.310 1405.200 1307.630 ;
        RECT 2297.800 1307.310 2298.060 1307.630 ;
        RECT 2297.860 17.410 2298.000 1307.310 ;
        RECT 2297.860 17.270 2298.460 17.410 ;
        RECT 2298.320 2.400 2298.460 17.270 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
      LAYER via2 ;
        RECT 1190.570 1335.040 1190.850 1335.320 ;
        RECT 1405.390 1335.040 1405.670 1335.320 ;
      LAYER met3 ;
        RECT 1190.545 1335.330 1190.875 1335.345 ;
        RECT 1405.365 1335.330 1405.695 1335.345 ;
        RECT 1190.545 1335.030 1405.695 1335.330 ;
        RECT 1190.545 1335.015 1190.875 1335.030 ;
        RECT 1405.365 1335.015 1405.695 1335.030 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1055.940 1421.330 1056.000 ;
        RECT 2311.570 1055.940 2311.890 1056.000 ;
        RECT 1421.010 1055.800 2311.890 1055.940 ;
        RECT 1421.010 1055.740 1421.330 1055.800 ;
        RECT 2311.570 1055.740 2311.890 1055.800 ;
      LAYER via ;
        RECT 1421.040 1055.740 1421.300 1056.000 ;
        RECT 2311.600 1055.740 2311.860 1056.000 ;
      LAYER met2 ;
        RECT 1421.030 1060.955 1421.310 1061.325 ;
        RECT 1421.100 1056.030 1421.240 1060.955 ;
        RECT 1421.040 1055.710 1421.300 1056.030 ;
        RECT 2311.600 1055.710 2311.860 1056.030 ;
        RECT 2311.660 17.410 2311.800 1055.710 ;
        RECT 2311.660 17.270 2316.400 17.410 ;
        RECT 2316.260 2.400 2316.400 17.270 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1061.000 1421.310 1061.280 ;
      LAYER met3 ;
        RECT 1421.005 1061.290 1421.335 1061.305 ;
        RECT 1408.060 1061.200 1421.335 1061.290 ;
        RECT 1404.305 1060.990 1421.335 1061.200 ;
        RECT 1404.305 1060.600 1408.305 1060.990 ;
        RECT 1421.005 1060.975 1421.335 1060.990 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 724.110 113.800 724.430 113.860 ;
        RECT 2332.270 113.800 2332.590 113.860 ;
        RECT 724.110 113.660 2332.590 113.800 ;
        RECT 724.110 113.600 724.430 113.660 ;
        RECT 2332.270 113.600 2332.590 113.660 ;
      LAYER via ;
        RECT 724.140 113.600 724.400 113.860 ;
        RECT 2332.300 113.600 2332.560 113.860 ;
      LAYER met2 ;
        RECT 723.170 216.650 723.450 220.000 ;
        RECT 723.170 216.510 724.340 216.650 ;
        RECT 723.170 216.000 723.450 216.510 ;
        RECT 724.200 113.890 724.340 216.510 ;
        RECT 724.140 113.570 724.400 113.890 ;
        RECT 2332.300 113.570 2332.560 113.890 ;
        RECT 2332.360 17.410 2332.500 113.570 ;
        RECT 2332.360 17.270 2334.340 17.410 ;
        RECT 2334.200 2.400 2334.340 17.270 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1420.090 448.700 1420.410 448.760 ;
        RECT 2346.070 448.700 2346.390 448.760 ;
        RECT 1420.090 448.560 2346.390 448.700 ;
        RECT 1420.090 448.500 1420.410 448.560 ;
        RECT 2346.070 448.500 2346.390 448.560 ;
      LAYER via ;
        RECT 1420.120 448.500 1420.380 448.760 ;
        RECT 2346.100 448.500 2346.360 448.760 ;
      LAYER met2 ;
        RECT 1420.110 454.395 1420.390 454.765 ;
        RECT 1420.180 448.790 1420.320 454.395 ;
        RECT 1420.120 448.470 1420.380 448.790 ;
        RECT 2346.100 448.470 2346.360 448.790 ;
        RECT 2346.160 17.410 2346.300 448.470 ;
        RECT 2346.160 17.270 2351.820 17.410 ;
        RECT 2351.680 2.400 2351.820 17.270 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
      LAYER via2 ;
        RECT 1420.110 454.440 1420.390 454.720 ;
      LAYER met3 ;
        RECT 1420.085 454.730 1420.415 454.745 ;
        RECT 1408.060 454.640 1420.415 454.730 ;
        RECT 1404.305 454.430 1420.415 454.640 ;
        RECT 1404.305 454.040 1408.305 454.430 ;
        RECT 1420.085 454.415 1420.415 454.430 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2366.790 127.995 2367.070 128.365 ;
        RECT 2366.860 17.410 2367.000 127.995 ;
        RECT 2366.860 17.270 2369.760 17.410 ;
        RECT 2369.620 2.400 2369.760 17.270 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
      LAYER via2 ;
        RECT 2366.790 128.040 2367.070 128.320 ;
      LAYER met3 ;
        RECT 310.000 241.880 314.000 242.480 ;
        RECT 311.270 241.220 311.570 241.880 ;
        RECT 311.230 240.900 311.610 241.220 ;
        RECT 311.230 219.450 311.610 219.460 ;
        RECT 314.910 219.450 315.290 219.460 ;
        RECT 311.230 219.150 315.290 219.450 ;
        RECT 311.230 219.140 311.610 219.150 ;
        RECT 314.910 219.140 315.290 219.150 ;
        RECT 314.910 128.330 315.290 128.340 ;
        RECT 2366.765 128.330 2367.095 128.345 ;
        RECT 314.910 128.030 2367.095 128.330 ;
        RECT 314.910 128.020 315.290 128.030 ;
        RECT 2366.765 128.015 2367.095 128.030 ;
      LAYER via3 ;
        RECT 311.260 240.900 311.580 241.220 ;
        RECT 311.260 219.140 311.580 219.460 ;
        RECT 314.940 219.140 315.260 219.460 ;
        RECT 314.940 128.020 315.260 128.340 ;
      LAYER met4 ;
        RECT 311.255 240.895 311.585 241.225 ;
        RECT 311.270 219.465 311.570 240.895 ;
        RECT 311.255 219.135 311.585 219.465 ;
        RECT 314.935 219.135 315.265 219.465 ;
        RECT 314.950 128.345 315.250 219.135 ;
        RECT 314.935 128.015 315.265 128.345 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 869.620 1421.330 869.680 ;
        RECT 2387.470 869.620 2387.790 869.680 ;
        RECT 1421.010 869.480 2387.790 869.620 ;
        RECT 1421.010 869.420 1421.330 869.480 ;
        RECT 2387.470 869.420 2387.790 869.480 ;
      LAYER via ;
        RECT 1421.040 869.420 1421.300 869.680 ;
        RECT 2387.500 869.420 2387.760 869.680 ;
      LAYER met2 ;
        RECT 1421.030 870.555 1421.310 870.925 ;
        RECT 1421.100 869.710 1421.240 870.555 ;
        RECT 1421.040 869.390 1421.300 869.710 ;
        RECT 2387.500 869.390 2387.760 869.710 ;
        RECT 2387.560 2.400 2387.700 869.390 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
      LAYER via2 ;
        RECT 1421.030 870.600 1421.310 870.880 ;
      LAYER met3 ;
        RECT 1421.005 870.890 1421.335 870.905 ;
        RECT 1408.060 870.800 1421.335 870.890 ;
        RECT 1404.305 870.590 1421.335 870.800 ;
        RECT 1404.305 870.200 1408.305 870.590 ;
        RECT 1421.005 870.575 1421.335 870.590 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2401.290 147.715 2401.570 148.085 ;
        RECT 2401.360 17.410 2401.500 147.715 ;
        RECT 2401.360 17.270 2405.640 17.410 ;
        RECT 2405.500 2.400 2405.640 17.270 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
      LAYER via2 ;
        RECT 2401.290 147.760 2401.570 148.040 ;
      LAYER met3 ;
        RECT 300.190 307.850 300.570 307.860 ;
        RECT 300.190 307.760 310.500 307.850 ;
        RECT 300.190 307.550 314.000 307.760 ;
        RECT 300.190 307.540 300.570 307.550 ;
        RECT 310.000 307.160 314.000 307.550 ;
        RECT 300.190 148.050 300.570 148.060 ;
        RECT 2401.265 148.050 2401.595 148.065 ;
        RECT 300.190 147.750 2401.595 148.050 ;
        RECT 300.190 147.740 300.570 147.750 ;
        RECT 2401.265 147.735 2401.595 147.750 ;
      LAYER via3 ;
        RECT 300.220 307.540 300.540 307.860 ;
        RECT 300.220 147.740 300.540 148.060 ;
      LAYER met4 ;
        RECT 300.215 307.535 300.545 307.865 ;
        RECT 300.230 148.065 300.530 307.535 ;
        RECT 300.215 147.735 300.545 148.065 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 799.550 39.680 799.870 39.740 ;
        RECT 1414.570 39.680 1414.890 39.740 ;
        RECT 799.550 39.540 1414.890 39.680 ;
        RECT 799.550 39.480 799.870 39.540 ;
        RECT 1414.570 39.480 1414.890 39.540 ;
      LAYER via ;
        RECT 799.580 39.480 799.840 39.740 ;
        RECT 1414.600 39.480 1414.860 39.740 ;
      LAYER met2 ;
        RECT 1414.590 1177.915 1414.870 1178.285 ;
        RECT 1414.660 39.770 1414.800 1177.915 ;
        RECT 799.580 39.450 799.840 39.770 ;
        RECT 1414.600 39.450 1414.860 39.770 ;
        RECT 799.640 2.400 799.780 39.450 ;
        RECT 799.430 -4.800 799.990 2.400 ;
      LAYER via2 ;
        RECT 1414.590 1177.960 1414.870 1178.240 ;
      LAYER met3 ;
        RECT 1414.565 1178.250 1414.895 1178.265 ;
        RECT 1408.060 1178.160 1414.895 1178.250 ;
        RECT 1404.305 1177.950 1414.895 1178.160 ;
        RECT 1404.305 1177.560 1408.305 1177.950 ;
        RECT 1414.565 1177.935 1414.895 1177.950 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 281.590 1334.060 281.910 1334.120 ;
        RECT 774.710 1334.060 775.030 1334.120 ;
        RECT 281.590 1333.920 775.030 1334.060 ;
        RECT 281.590 1333.860 281.910 1333.920 ;
        RECT 774.710 1333.860 775.030 1333.920 ;
        RECT 281.590 210.700 281.910 210.760 ;
        RECT 642.230 210.700 642.550 210.760 ;
        RECT 281.590 210.560 642.550 210.700 ;
        RECT 281.590 210.500 281.910 210.560 ;
        RECT 642.230 210.500 642.550 210.560 ;
        RECT 642.230 17.240 642.550 17.300 ;
        RECT 644.990 17.240 645.310 17.300 ;
        RECT 642.230 17.100 645.310 17.240 ;
        RECT 642.230 17.040 642.550 17.100 ;
        RECT 644.990 17.040 645.310 17.100 ;
      LAYER via ;
        RECT 281.620 1333.860 281.880 1334.120 ;
        RECT 774.740 1333.860 775.000 1334.120 ;
        RECT 281.620 210.500 281.880 210.760 ;
        RECT 642.260 210.500 642.520 210.760 ;
        RECT 642.260 17.040 642.520 17.300 ;
        RECT 645.020 17.040 645.280 17.300 ;
      LAYER met2 ;
        RECT 281.620 1333.830 281.880 1334.150 ;
        RECT 774.740 1333.830 775.000 1334.150 ;
        RECT 281.680 210.790 281.820 1333.830 ;
        RECT 774.800 1325.025 774.940 1333.830 ;
        RECT 774.690 1321.025 774.970 1325.025 ;
        RECT 281.620 210.470 281.880 210.790 ;
        RECT 642.260 210.470 642.520 210.790 ;
        RECT 642.320 17.330 642.460 210.470 ;
        RECT 642.260 17.010 642.520 17.330 ;
        RECT 645.020 17.010 645.280 17.330 ;
        RECT 645.080 2.400 645.220 17.010 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1406.290 1300.740 1406.610 1300.800 ;
        RECT 2428.870 1300.740 2429.190 1300.800 ;
        RECT 1406.290 1300.600 2429.190 1300.740 ;
        RECT 1406.290 1300.540 1406.610 1300.600 ;
        RECT 2428.870 1300.540 2429.190 1300.600 ;
      LAYER via ;
        RECT 1406.320 1300.540 1406.580 1300.800 ;
        RECT 2428.900 1300.540 2429.160 1300.800 ;
      LAYER met2 ;
        RECT 518.050 1333.635 518.330 1334.005 ;
        RECT 1406.310 1333.635 1406.590 1334.005 ;
        RECT 518.120 1325.025 518.260 1333.635 ;
        RECT 518.010 1321.025 518.290 1325.025 ;
        RECT 1406.380 1300.830 1406.520 1333.635 ;
        RECT 1406.320 1300.510 1406.580 1300.830 ;
        RECT 2428.900 1300.510 2429.160 1300.830 ;
        RECT 2428.960 2.400 2429.100 1300.510 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
      LAYER via2 ;
        RECT 518.050 1333.680 518.330 1333.960 ;
        RECT 1406.310 1333.680 1406.590 1333.960 ;
      LAYER met3 ;
        RECT 518.025 1333.970 518.355 1333.985 ;
        RECT 1406.285 1333.970 1406.615 1333.985 ;
        RECT 518.025 1333.670 1406.615 1333.970 ;
        RECT 518.025 1333.655 518.355 1333.670 ;
        RECT 1406.285 1333.655 1406.615 1333.670 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 294.930 93.060 295.250 93.120 ;
        RECT 2442.670 93.060 2442.990 93.120 ;
        RECT 294.930 92.920 2442.990 93.060 ;
        RECT 294.930 92.860 295.250 92.920 ;
        RECT 2442.670 92.860 2442.990 92.920 ;
      LAYER via ;
        RECT 294.960 92.860 295.220 93.120 ;
        RECT 2442.700 92.860 2442.960 93.120 ;
      LAYER met2 ;
        RECT 294.950 929.035 295.230 929.405 ;
        RECT 295.020 93.150 295.160 929.035 ;
        RECT 294.960 92.830 295.220 93.150 ;
        RECT 2442.700 92.830 2442.960 93.150 ;
        RECT 2442.760 17.410 2442.900 92.830 ;
        RECT 2442.760 17.270 2447.040 17.410 ;
        RECT 2446.900 2.400 2447.040 17.270 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
      LAYER via2 ;
        RECT 294.950 929.080 295.230 929.360 ;
      LAYER met3 ;
        RECT 294.925 929.370 295.255 929.385 ;
        RECT 294.925 929.280 310.500 929.370 ;
        RECT 294.925 929.070 314.000 929.280 ;
        RECT 294.925 929.055 295.255 929.070 ;
        RECT 310.000 928.680 314.000 929.070 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1148.765 1320.985 1148.935 1321.835 ;
      LAYER mcon ;
        RECT 1148.765 1321.665 1148.935 1321.835 ;
      LAYER met1 ;
        RECT 1051.630 1332.020 1051.950 1332.080 ;
        RECT 1131.210 1332.020 1131.530 1332.080 ;
        RECT 1051.630 1331.880 1131.530 1332.020 ;
        RECT 1051.630 1331.820 1051.950 1331.880 ;
        RECT 1131.210 1331.820 1131.530 1331.880 ;
        RECT 1131.210 1321.820 1131.530 1321.880 ;
        RECT 1148.705 1321.820 1148.995 1321.865 ;
        RECT 1131.210 1321.680 1148.995 1321.820 ;
        RECT 1131.210 1321.620 1131.530 1321.680 ;
        RECT 1148.705 1321.635 1148.995 1321.680 ;
        RECT 1148.705 1321.140 1148.995 1321.185 ;
        RECT 2463.370 1321.140 2463.690 1321.200 ;
        RECT 1148.705 1321.000 2463.690 1321.140 ;
        RECT 1148.705 1320.955 1148.995 1321.000 ;
        RECT 2463.370 1320.940 2463.690 1321.000 ;
      LAYER via ;
        RECT 1051.660 1331.820 1051.920 1332.080 ;
        RECT 1131.240 1331.820 1131.500 1332.080 ;
        RECT 1131.240 1321.620 1131.500 1321.880 ;
        RECT 2463.400 1320.940 2463.660 1321.200 ;
      LAYER met2 ;
        RECT 1051.660 1331.790 1051.920 1332.110 ;
        RECT 1131.240 1331.790 1131.500 1332.110 ;
        RECT 1051.720 1325.025 1051.860 1331.790 ;
        RECT 1051.610 1321.025 1051.890 1325.025 ;
        RECT 1131.300 1321.910 1131.440 1331.790 ;
        RECT 1131.240 1321.590 1131.500 1321.910 ;
        RECT 2463.400 1320.910 2463.660 1321.230 ;
        RECT 2463.460 16.730 2463.600 1320.910 ;
        RECT 2463.460 16.590 2464.980 16.730 ;
        RECT 2464.840 2.400 2464.980 16.590 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 779.310 1329.300 779.630 1329.360 ;
        RECT 2411.390 1329.300 2411.710 1329.360 ;
        RECT 779.310 1329.160 2411.710 1329.300 ;
        RECT 779.310 1329.100 779.630 1329.160 ;
        RECT 2411.390 1329.100 2411.710 1329.160 ;
        RECT 2411.850 17.240 2412.170 17.300 ;
        RECT 2482.690 17.240 2483.010 17.300 ;
        RECT 2411.850 17.100 2483.010 17.240 ;
        RECT 2411.850 17.040 2412.170 17.100 ;
        RECT 2482.690 17.040 2483.010 17.100 ;
      LAYER via ;
        RECT 779.340 1329.100 779.600 1329.360 ;
        RECT 2411.420 1329.100 2411.680 1329.360 ;
        RECT 2411.880 17.040 2412.140 17.300 ;
        RECT 2482.720 17.040 2482.980 17.300 ;
      LAYER met2 ;
        RECT 779.340 1329.070 779.600 1329.390 ;
        RECT 2411.420 1329.070 2411.680 1329.390 ;
        RECT 779.400 1325.025 779.540 1329.070 ;
        RECT 779.290 1321.025 779.570 1325.025 ;
        RECT 2411.480 25.570 2411.620 1329.070 ;
        RECT 2411.480 25.430 2412.080 25.570 ;
        RECT 2411.940 17.330 2412.080 25.430 ;
        RECT 2411.880 17.010 2412.140 17.330 ;
        RECT 2482.720 17.010 2482.980 17.330 ;
        RECT 2482.780 2.400 2482.920 17.010 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1358.985 1315.545 1359.155 1331.355 ;
      LAYER mcon ;
        RECT 1358.985 1331.185 1359.155 1331.355 ;
      LAYER met1 ;
        RECT 1358.910 1331.340 1359.230 1331.400 ;
        RECT 1358.715 1331.200 1359.230 1331.340 ;
        RECT 1358.910 1331.140 1359.230 1331.200 ;
        RECT 1358.925 1315.700 1359.215 1315.745 ;
        RECT 2497.870 1315.700 2498.190 1315.760 ;
        RECT 1358.925 1315.560 2498.190 1315.700 ;
        RECT 1358.925 1315.515 1359.215 1315.560 ;
        RECT 2497.870 1315.500 2498.190 1315.560 ;
      LAYER via ;
        RECT 1358.940 1331.140 1359.200 1331.400 ;
        RECT 2497.900 1315.500 2498.160 1315.760 ;
      LAYER met2 ;
        RECT 1289.010 1331.595 1289.290 1331.965 ;
        RECT 1358.930 1331.595 1359.210 1331.965 ;
        RECT 1289.080 1325.025 1289.220 1331.595 ;
        RECT 1359.000 1331.430 1359.140 1331.595 ;
        RECT 1358.940 1331.110 1359.200 1331.430 ;
        RECT 1288.970 1321.025 1289.250 1325.025 ;
        RECT 2497.900 1315.470 2498.160 1315.790 ;
        RECT 2497.960 17.410 2498.100 1315.470 ;
        RECT 2497.960 17.270 2500.860 17.410 ;
        RECT 2500.720 2.400 2500.860 17.270 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
      LAYER via2 ;
        RECT 1289.010 1331.640 1289.290 1331.920 ;
        RECT 1358.930 1331.640 1359.210 1331.920 ;
      LAYER met3 ;
        RECT 1288.985 1331.930 1289.315 1331.945 ;
        RECT 1358.905 1331.930 1359.235 1331.945 ;
        RECT 1288.985 1331.630 1359.235 1331.930 ;
        RECT 1288.985 1331.615 1289.315 1331.630 ;
        RECT 1358.905 1331.615 1359.235 1331.630 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 787.590 200.500 787.910 200.560 ;
        RECT 792.650 200.500 792.970 200.560 ;
        RECT 787.590 200.360 792.970 200.500 ;
        RECT 787.590 200.300 787.910 200.360 ;
        RECT 792.650 200.300 792.970 200.360 ;
        RECT 792.650 141.340 792.970 141.400 ;
        RECT 2512.130 141.340 2512.450 141.400 ;
        RECT 792.650 141.200 2512.450 141.340 ;
        RECT 792.650 141.140 792.970 141.200 ;
        RECT 2512.130 141.140 2512.450 141.200 ;
        RECT 2512.130 17.920 2512.450 17.980 ;
        RECT 2518.110 17.920 2518.430 17.980 ;
        RECT 2512.130 17.780 2518.430 17.920 ;
        RECT 2512.130 17.720 2512.450 17.780 ;
        RECT 2518.110 17.720 2518.430 17.780 ;
      LAYER via ;
        RECT 787.620 200.300 787.880 200.560 ;
        RECT 792.680 200.300 792.940 200.560 ;
        RECT 792.680 141.140 792.940 141.400 ;
        RECT 2512.160 141.140 2512.420 141.400 ;
        RECT 2512.160 17.720 2512.420 17.980 ;
        RECT 2518.140 17.720 2518.400 17.980 ;
      LAYER met2 ;
        RECT 787.570 216.000 787.850 220.000 ;
        RECT 787.680 200.590 787.820 216.000 ;
        RECT 787.620 200.270 787.880 200.590 ;
        RECT 792.680 200.270 792.940 200.590 ;
        RECT 792.740 141.430 792.880 200.270 ;
        RECT 792.680 141.110 792.940 141.430 ;
        RECT 2512.160 141.110 2512.420 141.430 ;
        RECT 2512.220 18.010 2512.360 141.110 ;
        RECT 2512.160 17.690 2512.420 18.010 ;
        RECT 2518.140 17.690 2518.400 18.010 ;
        RECT 2518.200 2.400 2518.340 17.690 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 220.900 1419.490 220.960 ;
        RECT 2532.370 220.900 2532.690 220.960 ;
        RECT 1419.170 220.760 2532.690 220.900 ;
        RECT 1419.170 220.700 1419.490 220.760 ;
        RECT 2532.370 220.700 2532.690 220.760 ;
      LAYER via ;
        RECT 1419.200 220.700 1419.460 220.960 ;
        RECT 2532.400 220.700 2532.660 220.960 ;
      LAYER met2 ;
        RECT 1419.190 227.275 1419.470 227.645 ;
        RECT 1419.260 220.990 1419.400 227.275 ;
        RECT 1419.200 220.670 1419.460 220.990 ;
        RECT 2532.400 220.670 2532.660 220.990 ;
        RECT 2532.460 17.410 2532.600 220.670 ;
        RECT 2532.460 17.270 2536.280 17.410 ;
        RECT 2536.140 2.400 2536.280 17.270 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
      LAYER via2 ;
        RECT 1419.190 227.320 1419.470 227.600 ;
      LAYER met3 ;
        RECT 1419.165 227.610 1419.495 227.625 ;
        RECT 1408.060 227.520 1419.495 227.610 ;
        RECT 1404.305 227.310 1419.495 227.520 ;
        RECT 1404.305 226.920 1408.305 227.310 ;
        RECT 1419.165 227.295 1419.495 227.310 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 979.870 200.500 980.190 200.560 ;
        RECT 985.850 200.500 986.170 200.560 ;
        RECT 979.870 200.360 986.170 200.500 ;
        RECT 979.870 200.300 980.190 200.360 ;
        RECT 985.850 200.300 986.170 200.360 ;
        RECT 985.850 79.460 986.170 79.520 ;
        RECT 2553.070 79.460 2553.390 79.520 ;
        RECT 985.850 79.320 2553.390 79.460 ;
        RECT 985.850 79.260 986.170 79.320 ;
        RECT 2553.070 79.260 2553.390 79.320 ;
      LAYER via ;
        RECT 979.900 200.300 980.160 200.560 ;
        RECT 985.880 200.300 986.140 200.560 ;
        RECT 985.880 79.260 986.140 79.520 ;
        RECT 2553.100 79.260 2553.360 79.520 ;
      LAYER met2 ;
        RECT 979.850 216.000 980.130 220.000 ;
        RECT 979.960 200.590 980.100 216.000 ;
        RECT 979.900 200.270 980.160 200.590 ;
        RECT 985.880 200.270 986.140 200.590 ;
        RECT 985.940 79.550 986.080 200.270 ;
        RECT 985.880 79.230 986.140 79.550 ;
        RECT 2553.100 79.230 2553.360 79.550 ;
        RECT 2553.160 17.410 2553.300 79.230 ;
        RECT 2553.160 17.270 2554.220 17.410 ;
        RECT 2554.080 2.400 2554.220 17.270 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.110 86.260 517.430 86.320 ;
        RECT 2566.870 86.260 2567.190 86.320 ;
        RECT 517.110 86.120 2567.190 86.260 ;
        RECT 517.110 86.060 517.430 86.120 ;
        RECT 2566.870 86.060 2567.190 86.120 ;
      LAYER via ;
        RECT 517.140 86.060 517.400 86.320 ;
        RECT 2566.900 86.060 2567.160 86.320 ;
      LAYER met2 ;
        RECT 515.250 216.650 515.530 220.000 ;
        RECT 515.250 216.510 517.340 216.650 ;
        RECT 515.250 216.000 515.530 216.510 ;
        RECT 517.200 86.350 517.340 216.510 ;
        RECT 517.140 86.030 517.400 86.350 ;
        RECT 2566.900 86.030 2567.160 86.350 ;
        RECT 2566.960 18.090 2567.100 86.030 ;
        RECT 2566.960 17.950 2572.160 18.090 ;
        RECT 2572.020 2.400 2572.160 17.950 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 966.180 1421.330 966.240 ;
        RECT 2587.570 966.180 2587.890 966.240 ;
        RECT 1421.010 966.040 2587.890 966.180 ;
        RECT 1421.010 965.980 1421.330 966.040 ;
        RECT 2587.570 965.980 2587.890 966.040 ;
      LAYER via ;
        RECT 1421.040 965.980 1421.300 966.240 ;
        RECT 2587.600 965.980 2587.860 966.240 ;
      LAYER met2 ;
        RECT 1421.030 972.555 1421.310 972.925 ;
        RECT 1421.100 966.270 1421.240 972.555 ;
        RECT 1421.040 965.950 1421.300 966.270 ;
        RECT 2587.600 965.950 2587.860 966.270 ;
        RECT 2587.660 17.410 2587.800 965.950 ;
        RECT 2587.660 17.270 2589.640 17.410 ;
        RECT 2589.500 2.400 2589.640 17.270 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
      LAYER via2 ;
        RECT 1421.030 972.600 1421.310 972.880 ;
      LAYER met3 ;
        RECT 1421.005 972.890 1421.335 972.905 ;
        RECT 1408.060 972.800 1421.335 972.890 ;
        RECT 1404.305 972.590 1421.335 972.800 ;
        RECT 1404.305 972.200 1408.305 972.590 ;
        RECT 1421.005 972.575 1421.335 972.590 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 288.950 1334.740 289.270 1334.800 ;
        RECT 641.310 1334.740 641.630 1334.800 ;
        RECT 288.950 1334.600 641.630 1334.740 ;
        RECT 288.950 1334.540 289.270 1334.600 ;
        RECT 641.310 1334.540 641.630 1334.600 ;
        RECT 288.950 20.300 289.270 20.360 ;
        RECT 823.470 20.300 823.790 20.360 ;
        RECT 288.950 20.160 823.790 20.300 ;
        RECT 288.950 20.100 289.270 20.160 ;
        RECT 823.470 20.100 823.790 20.160 ;
      LAYER via ;
        RECT 288.980 1334.540 289.240 1334.800 ;
        RECT 641.340 1334.540 641.600 1334.800 ;
        RECT 288.980 20.100 289.240 20.360 ;
        RECT 823.500 20.100 823.760 20.360 ;
      LAYER met2 ;
        RECT 288.980 1334.510 289.240 1334.830 ;
        RECT 641.340 1334.510 641.600 1334.830 ;
        RECT 289.040 20.390 289.180 1334.510 ;
        RECT 641.400 1325.025 641.540 1334.510 ;
        RECT 641.290 1321.025 641.570 1325.025 ;
        RECT 288.980 20.070 289.240 20.390 ;
        RECT 823.500 20.070 823.760 20.390 ;
        RECT 823.560 2.400 823.700 20.070 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.750 1349.700 602.070 1349.760 ;
        RECT 2601.370 1349.700 2601.690 1349.760 ;
        RECT 601.750 1349.560 2601.690 1349.700 ;
        RECT 601.750 1349.500 602.070 1349.560 ;
        RECT 2601.370 1349.500 2601.690 1349.560 ;
        RECT 2601.370 18.260 2601.690 18.320 ;
        RECT 2607.350 18.260 2607.670 18.320 ;
        RECT 2601.370 18.120 2607.670 18.260 ;
        RECT 2601.370 18.060 2601.690 18.120 ;
        RECT 2607.350 18.060 2607.670 18.120 ;
      LAYER via ;
        RECT 601.780 1349.500 602.040 1349.760 ;
        RECT 2601.400 1349.500 2601.660 1349.760 ;
        RECT 2601.400 18.060 2601.660 18.320 ;
        RECT 2607.380 18.060 2607.640 18.320 ;
      LAYER met2 ;
        RECT 601.780 1349.470 602.040 1349.790 ;
        RECT 2601.400 1349.470 2601.660 1349.790 ;
        RECT 601.840 1325.025 601.980 1349.470 ;
        RECT 601.730 1321.025 602.010 1325.025 ;
        RECT 2601.460 18.350 2601.600 1349.470 ;
        RECT 2601.400 18.030 2601.660 18.350 ;
        RECT 2607.380 18.030 2607.640 18.350 ;
        RECT 2607.440 2.400 2607.580 18.030 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2625.310 23.955 2625.590 24.325 ;
        RECT 2625.380 2.400 2625.520 23.955 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
      LAYER via2 ;
        RECT 2625.310 24.000 2625.590 24.280 ;
      LAYER met3 ;
        RECT 294.670 805.610 295.050 805.620 ;
        RECT 294.670 805.520 310.500 805.610 ;
        RECT 294.670 805.310 314.000 805.520 ;
        RECT 294.670 805.300 295.050 805.310 ;
        RECT 310.000 804.920 314.000 805.310 ;
        RECT 294.670 24.290 295.050 24.300 ;
        RECT 2625.285 24.290 2625.615 24.305 ;
        RECT 294.670 23.990 2625.615 24.290 ;
        RECT 294.670 23.980 295.050 23.990 ;
        RECT 2625.285 23.975 2625.615 23.990 ;
      LAYER via3 ;
        RECT 294.700 805.300 295.020 805.620 ;
        RECT 294.700 23.980 295.020 24.300 ;
      LAYER met4 ;
        RECT 294.695 805.295 295.025 805.625 ;
        RECT 294.710 24.305 295.010 805.295 ;
        RECT 294.695 23.975 295.025 24.305 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1326.155 399.650 1326.525 ;
        RECT 2642.790 1326.155 2643.070 1326.525 ;
        RECT 399.440 1325.025 399.580 1326.155 ;
        RECT 399.330 1321.025 399.610 1325.025 ;
        RECT 2642.860 17.410 2643.000 1326.155 ;
        RECT 2642.860 17.270 2643.460 17.410 ;
        RECT 2643.320 2.400 2643.460 17.270 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
      LAYER via2 ;
        RECT 399.370 1326.200 399.650 1326.480 ;
        RECT 2642.790 1326.200 2643.070 1326.480 ;
      LAYER met3 ;
        RECT 399.345 1326.490 399.675 1326.505 ;
        RECT 2642.765 1326.490 2643.095 1326.505 ;
        RECT 399.345 1326.190 2643.095 1326.490 ;
        RECT 399.345 1326.175 399.675 1326.190 ;
        RECT 2642.765 1326.175 2643.095 1326.190 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 800.545 1331.865 800.715 1332.715 ;
      LAYER mcon ;
        RECT 800.545 1332.545 800.715 1332.715 ;
      LAYER met1 ;
        RECT 789.430 1332.700 789.750 1332.760 ;
        RECT 800.485 1332.700 800.775 1332.745 ;
        RECT 789.430 1332.560 800.775 1332.700 ;
        RECT 789.430 1332.500 789.750 1332.560 ;
        RECT 800.485 1332.515 800.775 1332.560 ;
        RECT 800.485 1332.020 800.775 1332.065 ;
        RECT 817.030 1332.020 817.350 1332.080 ;
        RECT 800.485 1331.880 817.350 1332.020 ;
        RECT 800.485 1331.835 800.775 1331.880 ;
        RECT 817.030 1331.820 817.350 1331.880 ;
      LAYER via ;
        RECT 789.460 1332.500 789.720 1332.760 ;
        RECT 817.060 1331.820 817.320 1332.080 ;
      LAYER met2 ;
        RECT 789.460 1332.470 789.720 1332.790 ;
        RECT 789.520 1325.025 789.660 1332.470 ;
        RECT 817.060 1331.790 817.320 1332.110 ;
        RECT 789.410 1321.025 789.690 1325.025 ;
        RECT 817.120 1321.765 817.260 1331.790 ;
        RECT 817.050 1321.395 817.330 1321.765 ;
        RECT 2656.590 1320.715 2656.870 1321.085 ;
        RECT 2656.660 17.410 2656.800 1320.715 ;
        RECT 2656.660 17.270 2661.400 17.410 ;
        RECT 2661.260 2.400 2661.400 17.270 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
      LAYER via2 ;
        RECT 817.050 1321.440 817.330 1321.720 ;
        RECT 2656.590 1320.760 2656.870 1321.040 ;
      LAYER met3 ;
        RECT 817.025 1321.730 817.355 1321.745 ;
        RECT 817.025 1321.415 817.570 1321.730 ;
        RECT 817.270 1321.050 817.570 1321.415 ;
        RECT 2656.565 1321.050 2656.895 1321.065 ;
        RECT 817.270 1320.750 2656.895 1321.050 ;
        RECT 2656.565 1320.735 2656.895 1320.750 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1221.520 1421.330 1221.580 ;
        RECT 2677.270 1221.520 2677.590 1221.580 ;
        RECT 1421.010 1221.380 2677.590 1221.520 ;
        RECT 1421.010 1221.320 1421.330 1221.380 ;
        RECT 2677.270 1221.320 2677.590 1221.380 ;
      LAYER via ;
        RECT 1421.040 1221.320 1421.300 1221.580 ;
        RECT 2677.300 1221.320 2677.560 1221.580 ;
      LAYER met2 ;
        RECT 1421.030 1221.435 1421.310 1221.805 ;
        RECT 1421.040 1221.290 1421.300 1221.435 ;
        RECT 2677.300 1221.290 2677.560 1221.610 ;
        RECT 2677.360 17.410 2677.500 1221.290 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1221.480 1421.310 1221.760 ;
      LAYER met3 ;
        RECT 1421.005 1221.770 1421.335 1221.785 ;
        RECT 1408.060 1221.680 1421.335 1221.770 ;
        RECT 1404.305 1221.470 1421.335 1221.680 ;
        RECT 1404.305 1221.080 1408.305 1221.470 ;
        RECT 1421.005 1221.455 1421.335 1221.470 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1007.660 1421.330 1007.720 ;
        RECT 1686.890 1007.660 1687.210 1007.720 ;
        RECT 1421.010 1007.520 1687.210 1007.660 ;
        RECT 1421.010 1007.460 1421.330 1007.520 ;
        RECT 1686.890 1007.460 1687.210 1007.520 ;
        RECT 1686.890 258.640 1687.210 258.700 ;
        RECT 2691.070 258.640 2691.390 258.700 ;
        RECT 1686.890 258.500 2691.390 258.640 ;
        RECT 1686.890 258.440 1687.210 258.500 ;
        RECT 2691.070 258.440 2691.390 258.500 ;
      LAYER via ;
        RECT 1421.040 1007.460 1421.300 1007.720 ;
        RECT 1686.920 1007.460 1687.180 1007.720 ;
        RECT 1686.920 258.440 1687.180 258.700 ;
        RECT 2691.100 258.440 2691.360 258.700 ;
      LAYER met2 ;
        RECT 1421.030 1009.275 1421.310 1009.645 ;
        RECT 1421.100 1007.750 1421.240 1009.275 ;
        RECT 1421.040 1007.430 1421.300 1007.750 ;
        RECT 1686.920 1007.430 1687.180 1007.750 ;
        RECT 1686.980 258.730 1687.120 1007.430 ;
        RECT 1686.920 258.410 1687.180 258.730 ;
        RECT 2691.100 258.410 2691.360 258.730 ;
        RECT 2691.160 17.410 2691.300 258.410 ;
        RECT 2691.160 17.270 2696.820 17.410 ;
        RECT 2696.680 2.400 2696.820 17.270 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1009.320 1421.310 1009.600 ;
      LAYER met3 ;
        RECT 1421.005 1009.610 1421.335 1009.625 ;
        RECT 1408.060 1009.520 1421.335 1009.610 ;
        RECT 1404.305 1009.310 1421.335 1009.520 ;
        RECT 1404.305 1008.920 1408.305 1009.310 ;
        RECT 1421.005 1009.295 1421.335 1009.310 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 815.190 1343.240 815.510 1343.300 ;
        RECT 2712.230 1343.240 2712.550 1343.300 ;
        RECT 815.190 1343.100 2712.550 1343.240 ;
        RECT 815.190 1343.040 815.510 1343.100 ;
        RECT 2712.230 1343.040 2712.550 1343.100 ;
      LAYER via ;
        RECT 815.220 1343.040 815.480 1343.300 ;
        RECT 2712.260 1343.040 2712.520 1343.300 ;
      LAYER met2 ;
        RECT 815.220 1343.010 815.480 1343.330 ;
        RECT 2712.260 1343.010 2712.520 1343.330 ;
        RECT 815.280 1325.050 815.420 1343.010 ;
        RECT 814.430 1325.025 815.420 1325.050 ;
        RECT 814.250 1324.910 815.420 1325.025 ;
        RECT 814.250 1321.025 814.530 1324.910 ;
        RECT 2712.320 17.410 2712.460 1343.010 ;
        RECT 2712.320 17.270 2714.760 17.410 ;
        RECT 2714.620 2.400 2714.760 17.270 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1358.910 155.620 1359.230 155.680 ;
        RECT 2732.470 155.620 2732.790 155.680 ;
        RECT 1358.910 155.480 2732.790 155.620 ;
        RECT 1358.910 155.420 1359.230 155.480 ;
        RECT 2732.470 155.420 2732.790 155.480 ;
      LAYER via ;
        RECT 1358.940 155.420 1359.200 155.680 ;
        RECT 2732.500 155.420 2732.760 155.680 ;
      LAYER met2 ;
        RECT 1356.130 216.650 1356.410 220.000 ;
        RECT 1356.130 216.510 1359.140 216.650 ;
        RECT 1356.130 216.000 1356.410 216.510 ;
        RECT 1359.000 155.710 1359.140 216.510 ;
        RECT 1358.940 155.390 1359.200 155.710 ;
        RECT 2732.500 155.390 2732.760 155.710 ;
        RECT 2732.560 2.400 2732.700 155.390 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2746.270 2.960 2746.590 3.020 ;
        RECT 2750.410 2.960 2750.730 3.020 ;
        RECT 2746.270 2.820 2750.730 2.960 ;
        RECT 2746.270 2.760 2746.590 2.820 ;
        RECT 2750.410 2.760 2750.730 2.820 ;
      LAYER via ;
        RECT 2746.300 2.760 2746.560 3.020 ;
        RECT 2750.440 2.760 2750.700 3.020 ;
      LAYER met2 ;
        RECT 2746.290 79.035 2746.570 79.405 ;
        RECT 2746.360 3.050 2746.500 79.035 ;
        RECT 2746.300 2.730 2746.560 3.050 ;
        RECT 2750.440 2.730 2750.700 3.050 ;
        RECT 2750.500 2.400 2750.640 2.730 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
      LAYER via2 ;
        RECT 2746.290 79.080 2746.570 79.360 ;
      LAYER met3 ;
        RECT 292.830 724.010 293.210 724.020 ;
        RECT 292.830 723.920 310.500 724.010 ;
        RECT 292.830 723.710 314.000 723.920 ;
        RECT 292.830 723.700 293.210 723.710 ;
        RECT 310.000 723.320 314.000 723.710 ;
        RECT 292.830 79.370 293.210 79.380 ;
        RECT 2746.265 79.370 2746.595 79.385 ;
        RECT 292.830 79.070 2746.595 79.370 ;
        RECT 292.830 79.060 293.210 79.070 ;
        RECT 2746.265 79.055 2746.595 79.070 ;
      LAYER via3 ;
        RECT 292.860 723.700 293.180 724.020 ;
        RECT 292.860 79.060 293.180 79.380 ;
      LAYER met4 ;
        RECT 292.855 723.695 293.185 724.025 ;
        RECT 292.870 79.385 293.170 723.695 ;
        RECT 292.855 79.055 293.185 79.385 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 683.630 200.500 683.950 200.560 ;
        RECT 689.610 200.500 689.930 200.560 ;
        RECT 683.630 200.360 689.930 200.500 ;
        RECT 683.630 200.300 683.950 200.360 ;
        RECT 689.610 200.300 689.930 200.360 ;
        RECT 689.610 65.520 689.930 65.580 ;
        RECT 2766.970 65.520 2767.290 65.580 ;
        RECT 689.610 65.380 2767.290 65.520 ;
        RECT 689.610 65.320 689.930 65.380 ;
        RECT 2766.970 65.320 2767.290 65.380 ;
      LAYER via ;
        RECT 683.660 200.300 683.920 200.560 ;
        RECT 689.640 200.300 689.900 200.560 ;
        RECT 689.640 65.320 689.900 65.580 ;
        RECT 2767.000 65.320 2767.260 65.580 ;
      LAYER met2 ;
        RECT 683.610 216.000 683.890 220.000 ;
        RECT 683.720 200.590 683.860 216.000 ;
        RECT 683.660 200.270 683.920 200.590 ;
        RECT 689.640 200.270 689.900 200.590 ;
        RECT 689.700 65.610 689.840 200.270 ;
        RECT 689.640 65.290 689.900 65.610 ;
        RECT 2767.000 65.290 2767.260 65.610 ;
        RECT 2767.060 3.130 2767.200 65.290 ;
        RECT 2767.060 2.990 2768.120 3.130 ;
        RECT 2767.980 2.400 2768.120 2.990 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1076.470 1327.600 1076.790 1327.660 ;
        RECT 1430.670 1327.600 1430.990 1327.660 ;
        RECT 1076.470 1327.460 1430.990 1327.600 ;
        RECT 1076.470 1327.400 1076.790 1327.460 ;
        RECT 1430.670 1327.400 1430.990 1327.460 ;
        RECT 841.410 212.060 841.730 212.120 ;
        RECT 1430.670 212.060 1430.990 212.120 ;
        RECT 841.410 211.920 1430.990 212.060 ;
        RECT 841.410 211.860 841.730 211.920 ;
        RECT 1430.670 211.860 1430.990 211.920 ;
      LAYER via ;
        RECT 1076.500 1327.400 1076.760 1327.660 ;
        RECT 1430.700 1327.400 1430.960 1327.660 ;
        RECT 841.440 211.860 841.700 212.120 ;
        RECT 1430.700 211.860 1430.960 212.120 ;
      LAYER met2 ;
        RECT 1076.500 1327.370 1076.760 1327.690 ;
        RECT 1430.700 1327.370 1430.960 1327.690 ;
        RECT 1076.560 1325.025 1076.700 1327.370 ;
        RECT 1076.450 1321.025 1076.730 1325.025 ;
        RECT 1430.760 212.150 1430.900 1327.370 ;
        RECT 841.440 211.830 841.700 212.150 ;
        RECT 1430.700 211.830 1430.960 212.150 ;
        RECT 841.500 17.410 841.640 211.830 ;
        RECT 841.040 17.270 841.640 17.410 ;
        RECT 841.040 2.400 841.180 17.270 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1404.910 1316.040 1405.230 1316.100 ;
        RECT 2780.770 1316.040 2781.090 1316.100 ;
        RECT 1404.910 1315.900 2781.090 1316.040 ;
        RECT 1404.910 1315.840 1405.230 1315.900 ;
        RECT 2780.770 1315.840 2781.090 1315.900 ;
        RECT 2780.770 2.960 2781.090 3.020 ;
        RECT 2785.830 2.960 2786.150 3.020 ;
        RECT 2780.770 2.820 2786.150 2.960 ;
        RECT 2780.770 2.760 2781.090 2.820 ;
        RECT 2785.830 2.760 2786.150 2.820 ;
      LAYER via ;
        RECT 1404.940 1315.840 1405.200 1316.100 ;
        RECT 2780.800 1315.840 2781.060 1316.100 ;
        RECT 2780.800 2.760 2781.060 3.020 ;
        RECT 2785.860 2.760 2786.120 3.020 ;
      LAYER met2 ;
        RECT 1323.970 1336.355 1324.250 1336.725 ;
        RECT 1324.040 1325.025 1324.180 1336.355 ;
        RECT 1323.930 1321.025 1324.210 1325.025 ;
        RECT 1404.930 1317.315 1405.210 1317.685 ;
        RECT 1405.000 1316.130 1405.140 1317.315 ;
        RECT 1404.940 1315.810 1405.200 1316.130 ;
        RECT 2780.800 1315.810 2781.060 1316.130 ;
        RECT 2780.860 3.050 2781.000 1315.810 ;
        RECT 2780.800 2.730 2781.060 3.050 ;
        RECT 2785.860 2.730 2786.120 3.050 ;
        RECT 2785.920 2.400 2786.060 2.730 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
      LAYER via2 ;
        RECT 1323.970 1336.400 1324.250 1336.680 ;
        RECT 1404.930 1317.360 1405.210 1317.640 ;
      LAYER met3 ;
        RECT 1323.945 1336.690 1324.275 1336.705 ;
        RECT 1393.150 1336.690 1393.530 1336.700 ;
        RECT 1323.945 1336.390 1393.530 1336.690 ;
        RECT 1323.945 1336.375 1324.275 1336.390 ;
        RECT 1393.150 1336.380 1393.530 1336.390 ;
        RECT 1393.150 1317.650 1393.530 1317.660 ;
        RECT 1404.905 1317.650 1405.235 1317.665 ;
        RECT 1393.150 1317.350 1405.235 1317.650 ;
        RECT 1393.150 1317.340 1393.530 1317.350 ;
        RECT 1404.905 1317.335 1405.235 1317.350 ;
      LAYER via3 ;
        RECT 1393.180 1336.380 1393.500 1336.700 ;
        RECT 1393.180 1317.340 1393.500 1317.660 ;
      LAYER met4 ;
        RECT 1393.175 1336.375 1393.505 1336.705 ;
        RECT 1393.190 1317.665 1393.490 1336.375 ;
        RECT 1393.175 1317.335 1393.505 1317.665 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1418.250 496.980 1418.570 497.040 ;
        RECT 2770.190 496.980 2770.510 497.040 ;
        RECT 1418.250 496.840 2770.510 496.980 ;
        RECT 1418.250 496.780 1418.570 496.840 ;
        RECT 2770.190 496.780 2770.510 496.840 ;
        RECT 2770.190 65.520 2770.510 65.580 ;
        RECT 2801.470 65.520 2801.790 65.580 ;
        RECT 2770.190 65.380 2801.790 65.520 ;
        RECT 2770.190 65.320 2770.510 65.380 ;
        RECT 2801.470 65.320 2801.790 65.380 ;
      LAYER via ;
        RECT 1418.280 496.780 1418.540 497.040 ;
        RECT 2770.220 496.780 2770.480 497.040 ;
        RECT 2770.220 65.320 2770.480 65.580 ;
        RECT 2801.500 65.320 2801.760 65.580 ;
      LAYER met2 ;
        RECT 1418.270 497.915 1418.550 498.285 ;
        RECT 1418.340 497.070 1418.480 497.915 ;
        RECT 1418.280 496.750 1418.540 497.070 ;
        RECT 2770.220 496.750 2770.480 497.070 ;
        RECT 2770.280 65.610 2770.420 496.750 ;
        RECT 2770.220 65.290 2770.480 65.610 ;
        RECT 2801.500 65.290 2801.760 65.610 ;
        RECT 2801.560 17.410 2801.700 65.290 ;
        RECT 2801.560 17.270 2804.000 17.410 ;
        RECT 2803.860 2.400 2804.000 17.270 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
      LAYER via2 ;
        RECT 1418.270 497.960 1418.550 498.240 ;
      LAYER met3 ;
        RECT 1418.245 498.250 1418.575 498.265 ;
        RECT 1408.060 498.160 1418.575 498.250 ;
        RECT 1404.305 497.950 1418.575 498.160 ;
        RECT 1404.305 497.560 1408.305 497.950 ;
        RECT 1418.245 497.935 1418.575 497.950 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2815.730 17.920 2816.050 17.980 ;
        RECT 2821.710 17.920 2822.030 17.980 ;
        RECT 2815.730 17.780 2822.030 17.920 ;
        RECT 2815.730 17.720 2816.050 17.780 ;
        RECT 2821.710 17.720 2822.030 17.780 ;
      LAYER via ;
        RECT 2815.760 17.720 2816.020 17.980 ;
        RECT 2821.740 17.720 2822.000 17.980 ;
      LAYER met2 ;
        RECT 2815.750 120.515 2816.030 120.885 ;
        RECT 2815.820 18.010 2815.960 120.515 ;
        RECT 2815.760 17.690 2816.020 18.010 ;
        RECT 2821.740 17.690 2822.000 18.010 ;
        RECT 2821.800 2.400 2821.940 17.690 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
      LAYER via2 ;
        RECT 2815.750 120.560 2816.030 120.840 ;
      LAYER met3 ;
        RECT 293.750 855.930 294.130 855.940 ;
        RECT 293.750 855.840 310.500 855.930 ;
        RECT 293.750 855.630 314.000 855.840 ;
        RECT 293.750 855.620 294.130 855.630 ;
        RECT 310.000 855.240 314.000 855.630 ;
        RECT 293.750 120.850 294.130 120.860 ;
        RECT 2815.725 120.850 2816.055 120.865 ;
        RECT 293.750 120.550 2816.055 120.850 ;
        RECT 293.750 120.540 294.130 120.550 ;
        RECT 2815.725 120.535 2816.055 120.550 ;
      LAYER via3 ;
        RECT 293.780 855.620 294.100 855.940 ;
        RECT 293.780 120.540 294.100 120.860 ;
      LAYER met4 ;
        RECT 293.775 855.615 294.105 855.945 ;
        RECT 293.790 120.865 294.090 855.615 ;
        RECT 293.775 120.535 294.105 120.865 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 809.670 1325.900 809.990 1325.960 ;
        RECT 2176.790 1325.900 2177.110 1325.960 ;
        RECT 809.670 1325.760 2177.110 1325.900 ;
        RECT 809.670 1325.700 809.990 1325.760 ;
        RECT 2176.790 1325.700 2177.110 1325.760 ;
        RECT 2176.790 17.580 2177.110 17.640 ;
        RECT 2839.190 17.580 2839.510 17.640 ;
        RECT 2176.790 17.440 2839.510 17.580 ;
        RECT 2176.790 17.380 2177.110 17.440 ;
        RECT 2839.190 17.380 2839.510 17.440 ;
      LAYER via ;
        RECT 809.700 1325.700 809.960 1325.960 ;
        RECT 2176.820 1325.700 2177.080 1325.960 ;
        RECT 2176.820 17.380 2177.080 17.640 ;
        RECT 2839.220 17.380 2839.480 17.640 ;
      LAYER met2 ;
        RECT 809.700 1325.670 809.960 1325.990 ;
        RECT 2176.820 1325.670 2177.080 1325.990 ;
        RECT 809.760 1325.025 809.900 1325.670 ;
        RECT 809.650 1321.025 809.930 1325.025 ;
        RECT 2176.880 17.670 2177.020 1325.670 ;
        RECT 2176.820 17.350 2177.080 17.670 ;
        RECT 2839.220 17.350 2839.480 17.670 ;
        RECT 2839.280 2.400 2839.420 17.350 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2856.690 161.995 2856.970 162.365 ;
        RECT 2856.760 17.410 2856.900 161.995 ;
        RECT 2856.760 17.270 2857.360 17.410 ;
        RECT 2857.220 2.400 2857.360 17.270 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
      LAYER via2 ;
        RECT 2856.690 162.040 2856.970 162.320 ;
      LAYER met3 ;
        RECT 295.590 1002.810 295.970 1002.820 ;
        RECT 295.590 1002.720 310.500 1002.810 ;
        RECT 295.590 1002.510 314.000 1002.720 ;
        RECT 295.590 1002.500 295.970 1002.510 ;
        RECT 310.000 1002.120 314.000 1002.510 ;
        RECT 295.590 162.330 295.970 162.340 ;
        RECT 2856.665 162.330 2856.995 162.345 ;
        RECT 295.590 162.030 2856.995 162.330 ;
        RECT 295.590 162.020 295.970 162.030 ;
        RECT 2856.665 162.015 2856.995 162.030 ;
      LAYER via3 ;
        RECT 295.620 1002.500 295.940 1002.820 ;
        RECT 295.620 162.020 295.940 162.340 ;
      LAYER met4 ;
        RECT 295.615 1002.495 295.945 1002.825 ;
        RECT 295.630 162.345 295.930 1002.495 ;
        RECT 295.615 162.015 295.945 162.345 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1283.010 44.780 1283.330 44.840 ;
        RECT 2875.070 44.780 2875.390 44.840 ;
        RECT 1283.010 44.640 2875.390 44.780 ;
        RECT 1283.010 44.580 1283.330 44.640 ;
        RECT 2875.070 44.580 2875.390 44.640 ;
      LAYER via ;
        RECT 1283.040 44.580 1283.300 44.840 ;
        RECT 2875.100 44.580 2875.360 44.840 ;
      LAYER met2 ;
        RECT 1281.610 216.650 1281.890 220.000 ;
        RECT 1281.610 216.510 1283.240 216.650 ;
        RECT 1281.610 216.000 1281.890 216.510 ;
        RECT 1283.100 44.870 1283.240 216.510 ;
        RECT 1283.040 44.550 1283.300 44.870 ;
        RECT 2875.100 44.550 2875.360 44.870 ;
        RECT 2875.160 2.400 2875.300 44.550 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1398.930 1321.480 1399.250 1321.540 ;
        RECT 1403.990 1321.480 1404.310 1321.540 ;
        RECT 1398.930 1321.340 1404.310 1321.480 ;
        RECT 1398.930 1321.280 1399.250 1321.340 ;
        RECT 1403.990 1321.280 1404.310 1321.340 ;
        RECT 1403.990 1266.060 1404.310 1266.120 ;
        RECT 2891.170 1266.060 2891.490 1266.120 ;
        RECT 1403.990 1265.920 2891.490 1266.060 ;
        RECT 1403.990 1265.860 1404.310 1265.920 ;
        RECT 2891.170 1265.860 2891.490 1265.920 ;
      LAYER via ;
        RECT 1398.960 1321.280 1399.220 1321.540 ;
        RECT 1404.020 1321.280 1404.280 1321.540 ;
        RECT 1404.020 1265.860 1404.280 1266.120 ;
        RECT 2891.200 1265.860 2891.460 1266.120 ;
      LAYER met2 ;
        RECT 1397.530 1321.650 1397.810 1325.025 ;
        RECT 1397.530 1321.570 1399.160 1321.650 ;
        RECT 1397.530 1321.510 1399.220 1321.570 ;
        RECT 1397.530 1321.025 1397.810 1321.510 ;
        RECT 1398.960 1321.250 1399.220 1321.510 ;
        RECT 1404.020 1321.250 1404.280 1321.570 ;
        RECT 1404.080 1266.150 1404.220 1321.250 ;
        RECT 1404.020 1265.830 1404.280 1266.150 ;
        RECT 2891.200 1265.830 2891.460 1266.150 ;
        RECT 2891.260 3.130 2891.400 1265.830 ;
        RECT 2891.260 2.990 2893.240 3.130 ;
        RECT 2893.100 2.400 2893.240 2.990 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 359.790 1332.360 360.110 1332.420 ;
        RECT 1297.270 1332.360 1297.590 1332.420 ;
        RECT 359.790 1332.220 1297.590 1332.360 ;
        RECT 359.790 1332.160 360.110 1332.220 ;
        RECT 1297.270 1332.160 1297.590 1332.220 ;
        RECT 2905.430 2.960 2905.750 3.020 ;
        RECT 2910.950 2.960 2911.270 3.020 ;
        RECT 2905.430 2.820 2911.270 2.960 ;
        RECT 2905.430 2.760 2905.750 2.820 ;
        RECT 2910.950 2.760 2911.270 2.820 ;
      LAYER via ;
        RECT 359.820 1332.160 360.080 1332.420 ;
        RECT 1297.300 1332.160 1297.560 1332.420 ;
        RECT 2905.460 2.760 2905.720 3.020 ;
        RECT 2910.980 2.760 2911.240 3.020 ;
      LAYER met2 ;
        RECT 359.820 1332.130 360.080 1332.450 ;
        RECT 1297.300 1332.130 1297.560 1332.450 ;
        RECT 359.880 1325.025 360.020 1332.130 ;
        RECT 359.770 1321.025 360.050 1325.025 ;
        RECT 1297.360 1321.765 1297.500 1332.130 ;
        RECT 1341.450 1322.755 1341.730 1323.125 ;
        RECT 1399.410 1322.755 1399.690 1323.125 ;
        RECT 1341.520 1321.765 1341.660 1322.755 ;
        RECT 1399.480 1321.765 1399.620 1322.755 ;
        RECT 1297.290 1321.395 1297.570 1321.765 ;
        RECT 1341.450 1321.395 1341.730 1321.765 ;
        RECT 1399.410 1321.395 1399.690 1321.765 ;
        RECT 2905.450 1321.395 2905.730 1321.765 ;
        RECT 2905.520 3.050 2905.660 1321.395 ;
        RECT 2905.460 2.730 2905.720 3.050 ;
        RECT 2910.980 2.730 2911.240 3.050 ;
        RECT 2911.040 2.400 2911.180 2.730 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 1341.450 1322.800 1341.730 1323.080 ;
        RECT 1399.410 1322.800 1399.690 1323.080 ;
        RECT 1297.290 1321.440 1297.570 1321.720 ;
        RECT 1341.450 1321.440 1341.730 1321.720 ;
        RECT 1399.410 1321.440 1399.690 1321.720 ;
        RECT 2905.450 1321.440 2905.730 1321.720 ;
      LAYER met3 ;
        RECT 1341.425 1323.090 1341.755 1323.105 ;
        RECT 1399.385 1323.090 1399.715 1323.105 ;
        RECT 1341.425 1322.790 1399.715 1323.090 ;
        RECT 1341.425 1322.775 1341.755 1322.790 ;
        RECT 1399.385 1322.775 1399.715 1322.790 ;
        RECT 1297.265 1321.730 1297.595 1321.745 ;
        RECT 1341.425 1321.730 1341.755 1321.745 ;
        RECT 1297.265 1321.430 1341.755 1321.730 ;
        RECT 1297.265 1321.415 1297.595 1321.430 ;
        RECT 1341.425 1321.415 1341.755 1321.430 ;
        RECT 1399.385 1321.730 1399.715 1321.745 ;
        RECT 2905.425 1321.730 2905.755 1321.745 ;
        RECT 1399.385 1321.430 2905.755 1321.730 ;
        RECT 1399.385 1321.415 1399.715 1321.430 ;
        RECT 2905.425 1321.415 2905.755 1321.430 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 18.515 859.190 18.885 ;
        RECT 858.980 2.400 859.120 18.515 ;
        RECT 858.770 -4.800 859.330 2.400 ;
      LAYER via2 ;
        RECT 858.910 18.560 859.190 18.840 ;
      LAYER met3 ;
        RECT 298.350 1141.530 298.730 1141.540 ;
        RECT 298.350 1141.440 310.500 1141.530 ;
        RECT 298.350 1141.230 314.000 1141.440 ;
        RECT 298.350 1141.220 298.730 1141.230 ;
        RECT 310.000 1140.840 314.000 1141.230 ;
        RECT 320.430 159.610 320.810 159.620 ;
        RECT 320.430 159.310 321.690 159.610 ;
        RECT 320.430 159.300 320.810 159.310 ;
        RECT 321.390 158.940 321.690 159.310 ;
        RECT 321.350 158.620 321.730 158.940 ;
        RECT 321.350 96.740 321.730 97.060 ;
        RECT 321.390 95.700 321.690 96.740 ;
        RECT 321.350 95.380 321.730 95.700 ;
        RECT 319.510 18.850 319.890 18.860 ;
        RECT 858.885 18.850 859.215 18.865 ;
        RECT 319.510 18.550 859.215 18.850 ;
        RECT 319.510 18.540 319.890 18.550 ;
        RECT 858.885 18.535 859.215 18.550 ;
      LAYER via3 ;
        RECT 298.380 1141.220 298.700 1141.540 ;
        RECT 320.460 159.300 320.780 159.620 ;
        RECT 321.380 158.620 321.700 158.940 ;
        RECT 321.380 96.740 321.700 97.060 ;
        RECT 321.380 95.380 321.700 95.700 ;
        RECT 319.540 18.540 319.860 18.860 ;
      LAYER met4 ;
        RECT 298.375 1141.215 298.705 1141.545 ;
        RECT 298.390 342.290 298.690 1141.215 ;
        RECT 297.950 341.110 299.130 342.290 ;
        RECT 320.030 341.110 321.210 342.290 ;
        RECT 320.470 324.850 320.770 341.110 ;
        RECT 320.470 324.550 321.690 324.850 ;
        RECT 321.390 260.250 321.690 324.550 ;
        RECT 319.550 259.950 321.690 260.250 ;
        RECT 319.550 205.850 319.850 259.950 ;
        RECT 319.550 205.550 320.770 205.850 ;
        RECT 320.470 159.625 320.770 205.550 ;
        RECT 320.455 159.295 320.785 159.625 ;
        RECT 321.375 158.615 321.705 158.945 ;
        RECT 321.390 97.065 321.690 158.615 ;
        RECT 321.375 96.735 321.705 97.065 ;
        RECT 321.375 95.375 321.705 95.705 ;
        RECT 321.390 59.650 321.690 95.375 ;
        RECT 319.550 59.350 321.690 59.650 ;
        RECT 319.550 18.865 319.850 59.350 ;
        RECT 319.535 18.535 319.865 18.865 ;
      LAYER met5 ;
        RECT 297.740 340.900 321.420 342.500 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 882.810 115.160 883.130 115.220 ;
        RECT 1417.330 115.160 1417.650 115.220 ;
        RECT 882.810 115.020 1417.650 115.160 ;
        RECT 882.810 114.960 883.130 115.020 ;
        RECT 1417.330 114.960 1417.650 115.020 ;
        RECT 876.830 16.900 877.150 16.960 ;
        RECT 882.810 16.900 883.130 16.960 ;
        RECT 876.830 16.760 883.130 16.900 ;
        RECT 876.830 16.700 877.150 16.760 ;
        RECT 882.810 16.700 883.130 16.760 ;
      LAYER via ;
        RECT 882.840 114.960 883.100 115.220 ;
        RECT 1417.360 114.960 1417.620 115.220 ;
        RECT 876.860 16.700 877.120 16.960 ;
        RECT 882.840 16.700 883.100 16.960 ;
      LAYER met2 ;
        RECT 1417.350 636.635 1417.630 637.005 ;
        RECT 1417.420 115.250 1417.560 636.635 ;
        RECT 882.840 114.930 883.100 115.250 ;
        RECT 1417.360 114.930 1417.620 115.250 ;
        RECT 882.900 16.990 883.040 114.930 ;
        RECT 876.860 16.670 877.120 16.990 ;
        RECT 882.840 16.670 883.100 16.990 ;
        RECT 876.920 2.400 877.060 16.670 ;
        RECT 876.710 -4.800 877.270 2.400 ;
      LAYER via2 ;
        RECT 1417.350 636.680 1417.630 636.960 ;
      LAYER met3 ;
        RECT 1417.325 636.970 1417.655 636.985 ;
        RECT 1408.060 636.880 1417.655 636.970 ;
        RECT 1404.305 636.670 1417.655 636.880 ;
        RECT 1404.305 636.280 1408.305 636.670 ;
        RECT 1417.325 636.655 1417.655 636.670 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1404.525 628.405 1404.695 676.175 ;
        RECT 1404.525 593.045 1404.695 627.895 ;
        RECT 1404.525 531.505 1404.695 579.615 ;
        RECT 1404.525 483.225 1404.695 530.995 ;
        RECT 1404.985 448.205 1405.155 482.715 ;
        RECT 1404.525 386.325 1404.695 434.775 ;
        RECT 1404.985 338.385 1405.155 386.155 ;
        RECT 1404.525 303.025 1404.695 337.875 ;
      LAYER mcon ;
        RECT 1404.525 676.005 1404.695 676.175 ;
        RECT 1404.525 627.725 1404.695 627.895 ;
        RECT 1404.525 579.445 1404.695 579.615 ;
        RECT 1404.525 530.825 1404.695 530.995 ;
        RECT 1404.985 482.545 1405.155 482.715 ;
        RECT 1404.525 434.605 1404.695 434.775 ;
        RECT 1404.985 385.985 1405.155 386.155 ;
        RECT 1404.525 337.705 1404.695 337.875 ;
      LAYER met1 ;
        RECT 1404.465 676.160 1404.755 676.205 ;
        RECT 1404.910 676.160 1405.230 676.220 ;
        RECT 1404.465 676.020 1405.230 676.160 ;
        RECT 1404.465 675.975 1404.755 676.020 ;
        RECT 1404.910 675.960 1405.230 676.020 ;
        RECT 1404.450 628.560 1404.770 628.620 ;
        RECT 1404.255 628.420 1404.770 628.560 ;
        RECT 1404.450 628.360 1404.770 628.420 ;
        RECT 1404.450 627.880 1404.770 627.940 ;
        RECT 1404.255 627.740 1404.770 627.880 ;
        RECT 1404.450 627.680 1404.770 627.740 ;
        RECT 1404.450 593.200 1404.770 593.260 ;
        RECT 1404.255 593.060 1404.770 593.200 ;
        RECT 1404.450 593.000 1404.770 593.060 ;
        RECT 1404.465 579.600 1404.755 579.645 ;
        RECT 1404.910 579.600 1405.230 579.660 ;
        RECT 1404.465 579.460 1405.230 579.600 ;
        RECT 1404.465 579.415 1404.755 579.460 ;
        RECT 1404.910 579.400 1405.230 579.460 ;
        RECT 1404.450 531.660 1404.770 531.720 ;
        RECT 1404.255 531.520 1404.770 531.660 ;
        RECT 1404.450 531.460 1404.770 531.520 ;
        RECT 1404.450 530.980 1404.770 531.040 ;
        RECT 1404.255 530.840 1404.770 530.980 ;
        RECT 1404.450 530.780 1404.770 530.840 ;
        RECT 1404.465 483.380 1404.755 483.425 ;
        RECT 1404.910 483.380 1405.230 483.440 ;
        RECT 1404.465 483.240 1405.230 483.380 ;
        RECT 1404.465 483.195 1404.755 483.240 ;
        RECT 1404.910 483.180 1405.230 483.240 ;
        RECT 1404.910 482.700 1405.230 482.760 ;
        RECT 1404.715 482.560 1405.230 482.700 ;
        RECT 1404.910 482.500 1405.230 482.560 ;
        RECT 1404.910 448.360 1405.230 448.420 ;
        RECT 1404.715 448.220 1405.230 448.360 ;
        RECT 1404.910 448.160 1405.230 448.220 ;
        RECT 1404.465 434.760 1404.755 434.805 ;
        RECT 1404.910 434.760 1405.230 434.820 ;
        RECT 1404.465 434.620 1405.230 434.760 ;
        RECT 1404.465 434.575 1404.755 434.620 ;
        RECT 1404.910 434.560 1405.230 434.620 ;
        RECT 1404.450 386.480 1404.770 386.540 ;
        RECT 1404.255 386.340 1404.770 386.480 ;
        RECT 1404.450 386.280 1404.770 386.340 ;
        RECT 1404.910 386.140 1405.230 386.200 ;
        RECT 1404.715 386.000 1405.230 386.140 ;
        RECT 1404.910 385.940 1405.230 386.000 ;
        RECT 1404.450 338.540 1404.770 338.600 ;
        RECT 1404.925 338.540 1405.215 338.585 ;
        RECT 1404.450 338.400 1405.215 338.540 ;
        RECT 1404.450 338.340 1404.770 338.400 ;
        RECT 1404.925 338.355 1405.215 338.400 ;
        RECT 1404.450 337.860 1404.770 337.920 ;
        RECT 1404.255 337.720 1404.770 337.860 ;
        RECT 1404.450 337.660 1404.770 337.720 ;
        RECT 1404.465 303.180 1404.755 303.225 ;
        RECT 1404.910 303.180 1405.230 303.240 ;
        RECT 1404.465 303.040 1405.230 303.180 ;
        RECT 1404.465 302.995 1404.755 303.040 ;
        RECT 1404.910 302.980 1405.230 303.040 ;
        RECT 1404.910 255.240 1405.230 255.300 ;
        RECT 1406.750 255.240 1407.070 255.300 ;
        RECT 1404.910 255.100 1407.070 255.240 ;
        RECT 1404.910 255.040 1405.230 255.100 ;
        RECT 1406.750 255.040 1407.070 255.100 ;
        RECT 896.610 183.500 896.930 183.560 ;
        RECT 1407.210 183.500 1407.530 183.560 ;
        RECT 896.610 183.360 1407.530 183.500 ;
        RECT 896.610 183.300 896.930 183.360 ;
        RECT 1407.210 183.300 1407.530 183.360 ;
      LAYER via ;
        RECT 1404.940 675.960 1405.200 676.220 ;
        RECT 1404.480 628.360 1404.740 628.620 ;
        RECT 1404.480 627.680 1404.740 627.940 ;
        RECT 1404.480 593.000 1404.740 593.260 ;
        RECT 1404.940 579.400 1405.200 579.660 ;
        RECT 1404.480 531.460 1404.740 531.720 ;
        RECT 1404.480 530.780 1404.740 531.040 ;
        RECT 1404.940 483.180 1405.200 483.440 ;
        RECT 1404.940 482.500 1405.200 482.760 ;
        RECT 1404.940 448.160 1405.200 448.420 ;
        RECT 1404.940 434.560 1405.200 434.820 ;
        RECT 1404.480 386.280 1404.740 386.540 ;
        RECT 1404.940 385.940 1405.200 386.200 ;
        RECT 1404.480 338.340 1404.740 338.600 ;
        RECT 1404.480 337.660 1404.740 337.920 ;
        RECT 1404.940 302.980 1405.200 303.240 ;
        RECT 1404.940 255.040 1405.200 255.300 ;
        RECT 1406.780 255.040 1407.040 255.300 ;
        RECT 896.640 183.300 896.900 183.560 ;
        RECT 1407.240 183.300 1407.500 183.560 ;
      LAYER met2 ;
        RECT 1404.930 862.395 1405.210 862.765 ;
        RECT 1405.000 773.005 1405.140 862.395 ;
        RECT 1404.930 772.635 1405.210 773.005 ;
        RECT 1406.770 772.635 1407.050 773.005 ;
        RECT 1406.840 677.125 1406.980 772.635 ;
        RECT 1406.770 676.755 1407.050 677.125 ;
        RECT 1404.930 676.075 1405.210 676.445 ;
        RECT 1404.940 675.930 1405.200 676.075 ;
        RECT 1404.480 628.330 1404.740 628.650 ;
        RECT 1404.540 627.970 1404.680 628.330 ;
        RECT 1404.480 627.650 1404.740 627.970 ;
        RECT 1404.480 592.970 1404.740 593.290 ;
        RECT 1404.540 579.770 1404.680 592.970 ;
        RECT 1404.540 579.690 1405.140 579.770 ;
        RECT 1404.540 579.630 1405.200 579.690 ;
        RECT 1404.940 579.370 1405.200 579.630 ;
        RECT 1405.000 579.215 1405.140 579.370 ;
        RECT 1404.480 531.430 1404.740 531.750 ;
        RECT 1404.540 531.070 1404.680 531.430 ;
        RECT 1404.480 530.750 1404.740 531.070 ;
        RECT 1404.940 483.150 1405.200 483.470 ;
        RECT 1405.000 482.790 1405.140 483.150 ;
        RECT 1404.940 482.470 1405.200 482.790 ;
        RECT 1404.940 448.130 1405.200 448.450 ;
        RECT 1405.000 434.850 1405.140 448.130 ;
        RECT 1404.940 434.530 1405.200 434.850 ;
        RECT 1404.540 386.570 1405.140 386.650 ;
        RECT 1404.480 386.510 1405.140 386.570 ;
        RECT 1404.480 386.250 1404.740 386.510 ;
        RECT 1405.000 386.230 1405.140 386.510 ;
        RECT 1404.940 385.910 1405.200 386.230 ;
        RECT 1404.480 338.310 1404.740 338.630 ;
        RECT 1404.540 337.950 1404.680 338.310 ;
        RECT 1404.480 337.630 1404.740 337.950 ;
        RECT 1404.940 302.950 1405.200 303.270 ;
        RECT 1405.000 255.330 1405.140 302.950 ;
        RECT 1404.940 255.010 1405.200 255.330 ;
        RECT 1406.780 255.010 1407.040 255.330 ;
        RECT 1406.840 254.730 1406.980 255.010 ;
        RECT 1406.840 254.590 1407.440 254.730 ;
        RECT 1407.300 183.590 1407.440 254.590 ;
        RECT 896.640 183.270 896.900 183.590 ;
        RECT 1407.240 183.270 1407.500 183.590 ;
        RECT 896.700 17.410 896.840 183.270 ;
        RECT 894.860 17.270 896.840 17.410 ;
        RECT 894.860 2.400 895.000 17.270 ;
        RECT 894.650 -4.800 895.210 2.400 ;
      LAYER via2 ;
        RECT 1404.930 862.440 1405.210 862.720 ;
        RECT 1404.930 772.680 1405.210 772.960 ;
        RECT 1406.770 772.680 1407.050 772.960 ;
        RECT 1406.770 676.800 1407.050 677.080 ;
        RECT 1404.930 676.120 1405.210 676.400 ;
      LAYER met3 ;
        RECT 1404.305 863.400 1408.305 864.000 ;
        RECT 1405.150 862.745 1405.450 863.400 ;
        RECT 1404.905 862.430 1405.450 862.745 ;
        RECT 1404.905 862.415 1405.235 862.430 ;
        RECT 1404.905 772.970 1405.235 772.985 ;
        RECT 1406.745 772.970 1407.075 772.985 ;
        RECT 1404.905 772.670 1407.075 772.970 ;
        RECT 1404.905 772.655 1405.235 772.670 ;
        RECT 1406.745 772.655 1407.075 772.670 ;
        RECT 1406.745 677.090 1407.075 677.105 ;
        RECT 1405.150 676.790 1407.075 677.090 ;
        RECT 1405.150 676.425 1405.450 676.790 ;
        RECT 1406.745 676.775 1407.075 676.790 ;
        RECT 1404.905 676.110 1405.450 676.425 ;
        RECT 1404.905 676.095 1405.235 676.110 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 912.710 33.220 913.030 33.280 ;
        RECT 1228.270 33.220 1228.590 33.280 ;
        RECT 912.710 33.080 1228.590 33.220 ;
        RECT 912.710 33.020 913.030 33.080 ;
        RECT 1228.270 33.020 1228.590 33.080 ;
      LAYER via ;
        RECT 912.740 33.020 913.000 33.280 ;
        RECT 1228.300 33.020 1228.560 33.280 ;
      LAYER met2 ;
        RECT 1231.930 216.650 1232.210 220.000 ;
        RECT 1228.360 216.510 1232.210 216.650 ;
        RECT 1228.360 33.310 1228.500 216.510 ;
        RECT 1231.930 216.000 1232.210 216.510 ;
        RECT 912.740 32.990 913.000 33.310 ;
        RECT 1228.300 32.990 1228.560 33.310 ;
        RECT 912.800 2.400 912.940 32.990 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 289.410 1334.400 289.730 1334.460 ;
        RECT 685.470 1334.400 685.790 1334.460 ;
        RECT 289.410 1334.260 685.790 1334.400 ;
        RECT 289.410 1334.200 289.730 1334.260 ;
        RECT 685.470 1334.200 685.790 1334.260 ;
        RECT 289.410 19.620 289.730 19.680 ;
        RECT 930.190 19.620 930.510 19.680 ;
        RECT 289.410 19.480 930.510 19.620 ;
        RECT 289.410 19.420 289.730 19.480 ;
        RECT 930.190 19.420 930.510 19.480 ;
      LAYER via ;
        RECT 289.440 1334.200 289.700 1334.460 ;
        RECT 685.500 1334.200 685.760 1334.460 ;
        RECT 289.440 19.420 289.700 19.680 ;
        RECT 930.220 19.420 930.480 19.680 ;
      LAYER met2 ;
        RECT 289.440 1334.170 289.700 1334.490 ;
        RECT 685.500 1334.170 685.760 1334.490 ;
        RECT 289.500 19.710 289.640 1334.170 ;
        RECT 685.560 1325.025 685.700 1334.170 ;
        RECT 685.450 1321.025 685.730 1325.025 ;
        RECT 289.440 19.390 289.700 19.710 ;
        RECT 930.220 19.390 930.480 19.710 ;
        RECT 930.280 2.400 930.420 19.390 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 948.130 44.100 948.450 44.160 ;
        RECT 1207.570 44.100 1207.890 44.160 ;
        RECT 948.130 43.960 1207.890 44.100 ;
        RECT 948.130 43.900 948.450 43.960 ;
        RECT 1207.570 43.900 1207.890 43.960 ;
      LAYER via ;
        RECT 948.160 43.900 948.420 44.160 ;
        RECT 1207.600 43.900 1207.860 44.160 ;
      LAYER met2 ;
        RECT 1212.610 216.650 1212.890 220.000 ;
        RECT 1207.660 216.510 1212.890 216.650 ;
        RECT 1207.660 44.190 1207.800 216.510 ;
        RECT 1212.610 216.000 1212.890 216.510 ;
        RECT 948.160 43.870 948.420 44.190 ;
        RECT 1207.600 43.870 1207.860 44.190 ;
        RECT 948.220 2.400 948.360 43.870 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 972.510 14.180 972.830 14.240 ;
        RECT 966.160 14.040 972.830 14.180 ;
        RECT 966.160 13.900 966.300 14.040 ;
        RECT 972.510 13.980 972.830 14.040 ;
        RECT 966.070 13.640 966.390 13.900 ;
      LAYER via ;
        RECT 972.540 13.980 972.800 14.240 ;
        RECT 966.100 13.640 966.360 13.900 ;
      LAYER met2 ;
        RECT 1224.610 1347.235 1224.890 1347.605 ;
        RECT 1224.680 1325.025 1224.820 1347.235 ;
        RECT 1224.570 1321.025 1224.850 1325.025 ;
        RECT 972.530 196.675 972.810 197.045 ;
        RECT 972.600 14.270 972.740 196.675 ;
        RECT 972.540 13.950 972.800 14.270 ;
        RECT 966.100 13.610 966.360 13.930 ;
        RECT 966.160 2.400 966.300 13.610 ;
        RECT 965.950 -4.800 966.510 2.400 ;
      LAYER via2 ;
        RECT 1224.610 1347.280 1224.890 1347.560 ;
        RECT 972.530 196.720 972.810 197.000 ;
      LAYER met3 ;
        RECT 1224.585 1347.570 1224.915 1347.585 ;
        RECT 1394.070 1347.570 1394.450 1347.580 ;
        RECT 1224.585 1347.270 1394.450 1347.570 ;
        RECT 1224.585 1347.255 1224.915 1347.270 ;
        RECT 1394.070 1347.260 1394.450 1347.270 ;
        RECT 972.505 197.010 972.835 197.025 ;
        RECT 1394.070 197.010 1394.450 197.020 ;
        RECT 972.505 196.710 1394.450 197.010 ;
        RECT 972.505 196.695 972.835 196.710 ;
        RECT 1394.070 196.700 1394.450 196.710 ;
      LAYER via3 ;
        RECT 1394.100 1347.260 1394.420 1347.580 ;
        RECT 1394.100 196.700 1394.420 197.020 ;
      LAYER met4 ;
        RECT 1394.095 1347.255 1394.425 1347.585 ;
        RECT 1394.110 197.025 1394.410 1347.255 ;
        RECT 1394.095 196.695 1394.425 197.025 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 984.010 44.440 984.330 44.500 ;
        RECT 1255.870 44.440 1256.190 44.500 ;
        RECT 984.010 44.300 1256.190 44.440 ;
        RECT 984.010 44.240 984.330 44.300 ;
        RECT 1255.870 44.240 1256.190 44.300 ;
      LAYER via ;
        RECT 984.040 44.240 984.300 44.500 ;
        RECT 1255.900 44.240 1256.160 44.500 ;
      LAYER met2 ;
        RECT 1256.770 216.650 1257.050 220.000 ;
        RECT 1255.960 216.510 1257.050 216.650 ;
        RECT 1255.960 44.530 1256.100 216.510 ;
        RECT 1256.770 216.000 1257.050 216.510 ;
        RECT 984.040 44.210 984.300 44.530 ;
        RECT 1255.900 44.210 1256.160 44.530 ;
        RECT 984.100 2.400 984.240 44.210 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 496.025 48.365 496.195 137.955 ;
      LAYER mcon ;
        RECT 496.025 137.785 496.195 137.955 ;
      LAYER met1 ;
        RECT 495.030 186.560 495.350 186.620 ;
        RECT 496.410 186.560 496.730 186.620 ;
        RECT 495.030 186.420 496.730 186.560 ;
        RECT 495.030 186.360 495.350 186.420 ;
        RECT 496.410 186.360 496.730 186.420 ;
        RECT 495.965 137.940 496.255 137.985 ;
        RECT 496.410 137.940 496.730 138.000 ;
        RECT 495.965 137.800 496.730 137.940 ;
        RECT 495.965 137.755 496.255 137.800 ;
        RECT 496.410 137.740 496.730 137.800 ;
        RECT 495.950 48.520 496.270 48.580 ;
        RECT 495.755 48.380 496.270 48.520 ;
        RECT 495.950 48.320 496.270 48.380 ;
        RECT 568.260 15.400 614.400 15.540 ;
        RECT 495.950 15.200 496.270 15.260 ;
        RECT 568.260 15.200 568.400 15.400 ;
        RECT 495.950 15.060 568.400 15.200 ;
        RECT 614.260 15.200 614.400 15.400 ;
        RECT 662.930 15.200 663.250 15.260 ;
        RECT 614.260 15.060 663.250 15.200 ;
        RECT 495.950 15.000 496.270 15.060 ;
        RECT 662.930 15.000 663.250 15.060 ;
      LAYER via ;
        RECT 495.060 186.360 495.320 186.620 ;
        RECT 496.440 186.360 496.700 186.620 ;
        RECT 496.440 137.740 496.700 138.000 ;
        RECT 495.980 48.320 496.240 48.580 ;
        RECT 495.980 15.000 496.240 15.260 ;
        RECT 662.960 15.000 663.220 15.260 ;
      LAYER met2 ;
        RECT 495.010 216.000 495.290 220.000 ;
        RECT 495.120 186.650 495.260 216.000 ;
        RECT 495.060 186.330 495.320 186.650 ;
        RECT 496.440 186.330 496.700 186.650 ;
        RECT 496.500 138.030 496.640 186.330 ;
        RECT 496.440 137.710 496.700 138.030 ;
        RECT 495.980 48.290 496.240 48.610 ;
        RECT 496.040 15.290 496.180 48.290 ;
        RECT 495.980 14.970 496.240 15.290 ;
        RECT 662.960 14.970 663.220 15.290 ;
        RECT 663.020 2.400 663.160 14.970 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 1332.275 533.050 1332.645 ;
        RECT 532.840 1325.025 532.980 1332.275 ;
        RECT 532.730 1321.025 533.010 1325.025 ;
        RECT 1001.970 17.835 1002.250 18.205 ;
        RECT 1002.040 2.400 1002.180 17.835 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
      LAYER via2 ;
        RECT 532.770 1332.320 533.050 1332.600 ;
        RECT 1001.970 17.880 1002.250 18.160 ;
      LAYER met3 ;
        RECT 323.190 1332.610 323.570 1332.620 ;
        RECT 532.745 1332.610 533.075 1332.625 ;
        RECT 323.190 1332.310 533.075 1332.610 ;
        RECT 323.190 1332.300 323.570 1332.310 ;
        RECT 532.745 1332.295 533.075 1332.310 ;
        RECT 323.190 18.170 323.570 18.180 ;
        RECT 1001.945 18.170 1002.275 18.185 ;
        RECT 323.190 17.870 1002.275 18.170 ;
        RECT 323.190 17.860 323.570 17.870 ;
        RECT 1001.945 17.855 1002.275 17.870 ;
      LAYER via3 ;
        RECT 323.220 1332.300 323.540 1332.620 ;
        RECT 323.220 17.860 323.540 18.180 ;
      LAYER met4 ;
        RECT 323.215 1332.295 323.545 1332.625 ;
        RECT 323.230 18.185 323.530 1332.295 ;
        RECT 323.215 17.855 323.545 18.185 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1404.065 1000.705 1404.235 1048.815 ;
        RECT 1404.985 954.125 1405.155 1000.195 ;
        RECT 1404.525 241.485 1404.695 263.755 ;
      LAYER mcon ;
        RECT 1404.065 1048.645 1404.235 1048.815 ;
        RECT 1404.985 1000.025 1405.155 1000.195 ;
        RECT 1404.525 263.585 1404.695 263.755 ;
      LAYER met1 ;
        RECT 1404.450 1049.140 1404.770 1049.200 ;
        RECT 1405.830 1049.140 1406.150 1049.200 ;
        RECT 1404.450 1049.000 1406.150 1049.140 ;
        RECT 1404.450 1048.940 1404.770 1049.000 ;
        RECT 1405.830 1048.940 1406.150 1049.000 ;
        RECT 1403.990 1048.800 1404.310 1048.860 ;
        RECT 1403.795 1048.660 1404.310 1048.800 ;
        RECT 1403.990 1048.600 1404.310 1048.660 ;
        RECT 1404.005 1000.860 1404.295 1000.905 ;
        RECT 1404.910 1000.860 1405.230 1000.920 ;
        RECT 1404.005 1000.720 1405.230 1000.860 ;
        RECT 1404.005 1000.675 1404.295 1000.720 ;
        RECT 1404.910 1000.660 1405.230 1000.720 ;
        RECT 1404.910 1000.180 1405.230 1000.240 ;
        RECT 1404.715 1000.040 1405.230 1000.180 ;
        RECT 1404.910 999.980 1405.230 1000.040 ;
        RECT 1404.910 954.280 1405.230 954.340 ;
        RECT 1404.715 954.140 1405.230 954.280 ;
        RECT 1404.910 954.080 1405.230 954.140 ;
        RECT 1404.910 896.820 1405.230 896.880 ;
        RECT 1407.210 896.820 1407.530 896.880 ;
        RECT 1404.910 896.680 1407.530 896.820 ;
        RECT 1404.910 896.620 1405.230 896.680 ;
        RECT 1407.210 896.620 1407.530 896.680 ;
        RECT 1406.290 834.600 1406.610 834.660 ;
        RECT 1407.210 834.600 1407.530 834.660 ;
        RECT 1406.290 834.460 1407.530 834.600 ;
        RECT 1406.290 834.400 1406.610 834.460 ;
        RECT 1407.210 834.400 1407.530 834.460 ;
        RECT 1403.990 763.200 1404.310 763.260 ;
        RECT 1405.830 763.200 1406.150 763.260 ;
        RECT 1403.990 763.060 1406.150 763.200 ;
        RECT 1403.990 763.000 1404.310 763.060 ;
        RECT 1405.830 763.000 1406.150 763.060 ;
        RECT 1403.990 600.680 1404.310 600.740 ;
        RECT 1405.830 600.680 1406.150 600.740 ;
        RECT 1403.990 600.540 1406.150 600.680 ;
        RECT 1403.990 600.480 1404.310 600.540 ;
        RECT 1405.830 600.480 1406.150 600.540 ;
        RECT 1403.990 569.740 1404.310 569.800 ;
        RECT 1405.830 569.740 1406.150 569.800 ;
        RECT 1403.990 569.600 1406.150 569.740 ;
        RECT 1403.990 569.540 1404.310 569.600 ;
        RECT 1405.830 569.540 1406.150 569.600 ;
        RECT 1403.990 531.320 1404.310 531.380 ;
        RECT 1405.830 531.320 1406.150 531.380 ;
        RECT 1403.990 531.180 1406.150 531.320 ;
        RECT 1403.990 531.120 1404.310 531.180 ;
        RECT 1405.830 531.120 1406.150 531.180 ;
        RECT 1403.990 473.180 1404.310 473.240 ;
        RECT 1405.830 473.180 1406.150 473.240 ;
        RECT 1403.990 473.040 1406.150 473.180 ;
        RECT 1403.990 472.980 1404.310 473.040 ;
        RECT 1405.830 472.980 1406.150 473.040 ;
        RECT 1403.990 424.560 1404.310 424.620 ;
        RECT 1406.750 424.560 1407.070 424.620 ;
        RECT 1403.990 424.420 1407.070 424.560 ;
        RECT 1403.990 424.360 1404.310 424.420 ;
        RECT 1406.750 424.360 1407.070 424.420 ;
        RECT 1403.990 376.620 1404.310 376.680 ;
        RECT 1406.750 376.620 1407.070 376.680 ;
        RECT 1403.990 376.480 1407.070 376.620 ;
        RECT 1403.990 376.420 1404.310 376.480 ;
        RECT 1406.750 376.420 1407.070 376.480 ;
        RECT 1403.990 327.320 1404.310 327.380 ;
        RECT 1406.750 327.320 1407.070 327.380 ;
        RECT 1403.990 327.180 1407.070 327.320 ;
        RECT 1403.990 327.120 1404.310 327.180 ;
        RECT 1406.750 327.120 1407.070 327.180 ;
        RECT 1404.465 263.740 1404.755 263.785 ;
        RECT 1406.750 263.740 1407.070 263.800 ;
        RECT 1404.465 263.600 1407.070 263.740 ;
        RECT 1404.465 263.555 1404.755 263.600 ;
        RECT 1406.750 263.540 1407.070 263.600 ;
        RECT 1404.450 241.640 1404.770 241.700 ;
        RECT 1404.255 241.500 1404.770 241.640 ;
        RECT 1404.450 241.440 1404.770 241.500 ;
        RECT 1019.890 100.200 1020.210 100.260 ;
        RECT 1403.070 100.200 1403.390 100.260 ;
        RECT 1019.890 100.060 1403.390 100.200 ;
        RECT 1019.890 100.000 1020.210 100.060 ;
        RECT 1403.070 100.000 1403.390 100.060 ;
      LAYER via ;
        RECT 1404.480 1048.940 1404.740 1049.200 ;
        RECT 1405.860 1048.940 1406.120 1049.200 ;
        RECT 1404.020 1048.600 1404.280 1048.860 ;
        RECT 1404.940 1000.660 1405.200 1000.920 ;
        RECT 1404.940 999.980 1405.200 1000.240 ;
        RECT 1404.940 954.080 1405.200 954.340 ;
        RECT 1404.940 896.620 1405.200 896.880 ;
        RECT 1407.240 896.620 1407.500 896.880 ;
        RECT 1406.320 834.400 1406.580 834.660 ;
        RECT 1407.240 834.400 1407.500 834.660 ;
        RECT 1404.020 763.000 1404.280 763.260 ;
        RECT 1405.860 763.000 1406.120 763.260 ;
        RECT 1404.020 600.480 1404.280 600.740 ;
        RECT 1405.860 600.480 1406.120 600.740 ;
        RECT 1404.020 569.540 1404.280 569.800 ;
        RECT 1405.860 569.540 1406.120 569.800 ;
        RECT 1404.020 531.120 1404.280 531.380 ;
        RECT 1405.860 531.120 1406.120 531.380 ;
        RECT 1404.020 472.980 1404.280 473.240 ;
        RECT 1405.860 472.980 1406.120 473.240 ;
        RECT 1404.020 424.360 1404.280 424.620 ;
        RECT 1406.780 424.360 1407.040 424.620 ;
        RECT 1404.020 376.420 1404.280 376.680 ;
        RECT 1406.780 376.420 1407.040 376.680 ;
        RECT 1404.020 327.120 1404.280 327.380 ;
        RECT 1406.780 327.120 1407.040 327.380 ;
        RECT 1406.780 263.540 1407.040 263.800 ;
        RECT 1404.480 241.440 1404.740 241.700 ;
        RECT 1019.920 100.000 1020.180 100.260 ;
        RECT 1403.100 100.000 1403.360 100.260 ;
      LAYER met2 ;
        RECT 1405.850 1096.315 1406.130 1096.685 ;
        RECT 1405.920 1049.230 1406.060 1096.315 ;
        RECT 1404.480 1048.970 1404.740 1049.230 ;
        RECT 1404.080 1048.910 1404.740 1048.970 ;
        RECT 1405.860 1048.910 1406.120 1049.230 ;
        RECT 1404.080 1048.890 1404.680 1048.910 ;
        RECT 1404.020 1048.830 1404.680 1048.890 ;
        RECT 1404.020 1048.570 1404.280 1048.830 ;
        RECT 1404.080 1048.415 1404.220 1048.570 ;
        RECT 1404.940 1000.630 1405.200 1000.950 ;
        RECT 1405.000 1000.270 1405.140 1000.630 ;
        RECT 1404.940 999.950 1405.200 1000.270 ;
        RECT 1404.940 954.050 1405.200 954.370 ;
        RECT 1405.000 896.910 1405.140 954.050 ;
        RECT 1404.940 896.590 1405.200 896.910 ;
        RECT 1407.240 896.590 1407.500 896.910 ;
        RECT 1407.300 834.690 1407.440 896.590 ;
        RECT 1406.320 834.370 1406.580 834.690 ;
        RECT 1407.240 834.370 1407.500 834.690 ;
        RECT 1406.380 811.650 1406.520 834.370 ;
        RECT 1405.920 811.510 1406.520 811.650 ;
        RECT 1405.920 763.290 1406.060 811.510 ;
        RECT 1404.020 762.970 1404.280 763.290 ;
        RECT 1405.860 762.970 1406.120 763.290 ;
        RECT 1404.080 762.690 1404.220 762.970 ;
        RECT 1403.620 762.550 1404.220 762.690 ;
        RECT 1403.620 600.680 1403.760 762.550 ;
        RECT 1404.020 600.680 1404.280 600.770 ;
        RECT 1403.620 600.540 1404.280 600.680 ;
        RECT 1404.020 600.450 1404.280 600.540 ;
        RECT 1405.860 600.450 1406.120 600.770 ;
        RECT 1405.920 569.830 1406.060 600.450 ;
        RECT 1404.020 569.570 1404.280 569.830 ;
        RECT 1403.620 569.510 1404.280 569.570 ;
        RECT 1405.860 569.510 1406.120 569.830 ;
        RECT 1403.620 569.430 1404.220 569.510 ;
        RECT 1403.620 532.170 1403.760 569.430 ;
        RECT 1403.620 532.030 1404.220 532.170 ;
        RECT 1404.080 531.410 1404.220 532.030 ;
        RECT 1404.020 531.090 1404.280 531.410 ;
        RECT 1405.860 531.090 1406.120 531.410 ;
        RECT 1405.920 473.270 1406.060 531.090 ;
        RECT 1404.020 473.010 1404.280 473.270 ;
        RECT 1403.620 472.950 1404.280 473.010 ;
        RECT 1405.860 472.950 1406.120 473.270 ;
        RECT 1403.620 472.870 1404.220 472.950 ;
        RECT 1403.620 424.730 1403.760 472.870 ;
        RECT 1403.620 424.650 1404.220 424.730 ;
        RECT 1403.620 424.590 1404.280 424.650 ;
        RECT 1404.020 424.330 1404.280 424.590 ;
        RECT 1406.780 424.330 1407.040 424.650 ;
        RECT 1406.840 376.710 1406.980 424.330 ;
        RECT 1404.020 376.450 1404.280 376.710 ;
        RECT 1403.620 376.390 1404.280 376.450 ;
        RECT 1406.780 376.390 1407.040 376.710 ;
        RECT 1403.620 376.310 1404.220 376.390 ;
        RECT 1403.620 327.490 1403.760 376.310 ;
        RECT 1403.620 327.410 1404.220 327.490 ;
        RECT 1403.620 327.350 1404.280 327.410 ;
        RECT 1404.020 327.090 1404.280 327.350 ;
        RECT 1406.780 327.090 1407.040 327.410 ;
        RECT 1406.840 263.830 1406.980 327.090 ;
        RECT 1406.780 263.510 1407.040 263.830 ;
        RECT 1404.480 241.410 1404.740 241.730 ;
        RECT 1404.540 220.050 1404.680 241.410 ;
        RECT 1403.620 219.910 1404.680 220.050 ;
        RECT 1403.620 217.330 1403.760 219.910 ;
        RECT 1403.160 217.190 1403.760 217.330 ;
        RECT 1403.160 100.290 1403.300 217.190 ;
        RECT 1019.920 99.970 1020.180 100.290 ;
        RECT 1403.100 99.970 1403.360 100.290 ;
        RECT 1019.980 17.410 1020.120 99.970 ;
        RECT 1019.520 17.270 1020.120 17.410 ;
        RECT 1019.520 2.400 1019.660 17.270 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
      LAYER via2 ;
        RECT 1405.850 1096.360 1406.130 1096.640 ;
      LAYER met3 ;
        RECT 1404.305 1097.320 1408.305 1097.920 ;
        RECT 1405.150 1096.650 1405.450 1097.320 ;
        RECT 1405.825 1096.650 1406.155 1096.665 ;
        RECT 1405.150 1096.350 1406.155 1096.650 ;
        RECT 1405.825 1096.335 1406.155 1096.350 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1041.510 205.940 1041.830 206.000 ;
        RECT 1058.990 205.940 1059.310 206.000 ;
        RECT 1041.510 205.800 1059.310 205.940 ;
        RECT 1041.510 205.740 1041.830 205.800 ;
        RECT 1058.990 205.740 1059.310 205.800 ;
        RECT 1037.370 15.200 1037.690 15.260 ;
        RECT 1041.510 15.200 1041.830 15.260 ;
        RECT 1037.370 15.060 1041.830 15.200 ;
        RECT 1037.370 15.000 1037.690 15.060 ;
        RECT 1041.510 15.000 1041.830 15.060 ;
      LAYER via ;
        RECT 1041.540 205.740 1041.800 206.000 ;
        RECT 1059.020 205.740 1059.280 206.000 ;
        RECT 1037.400 15.000 1037.660 15.260 ;
        RECT 1041.540 15.000 1041.800 15.260 ;
      LAYER met2 ;
        RECT 1058.970 216.000 1059.250 220.000 ;
        RECT 1059.080 206.030 1059.220 216.000 ;
        RECT 1041.540 205.710 1041.800 206.030 ;
        RECT 1059.020 205.710 1059.280 206.030 ;
        RECT 1041.600 15.290 1041.740 205.710 ;
        RECT 1037.400 14.970 1037.660 15.290 ;
        RECT 1041.540 14.970 1041.800 15.290 ;
        RECT 1037.460 2.400 1037.600 14.970 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1055.310 218.520 1055.630 218.580 ;
        RECT 1415.490 218.520 1415.810 218.580 ;
        RECT 1055.310 218.380 1415.810 218.520 ;
        RECT 1055.310 218.320 1055.630 218.380 ;
        RECT 1415.490 218.320 1415.810 218.380 ;
      LAYER via ;
        RECT 1055.340 218.320 1055.600 218.580 ;
        RECT 1415.520 218.320 1415.780 218.580 ;
      LAYER met2 ;
        RECT 1415.510 1264.955 1415.790 1265.325 ;
        RECT 1415.580 218.610 1415.720 1264.955 ;
        RECT 1055.340 218.290 1055.600 218.610 ;
        RECT 1415.520 218.290 1415.780 218.610 ;
        RECT 1055.400 2.400 1055.540 218.290 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
      LAYER via2 ;
        RECT 1415.510 1265.000 1415.790 1265.280 ;
      LAYER met3 ;
        RECT 1415.485 1265.290 1415.815 1265.305 ;
        RECT 1408.060 1265.200 1415.815 1265.290 ;
        RECT 1404.305 1264.990 1415.815 1265.200 ;
        RECT 1404.305 1264.600 1408.305 1264.990 ;
        RECT 1415.485 1264.975 1415.815 1264.990 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1041.050 40.020 1041.370 40.080 ;
        RECT 1073.250 40.020 1073.570 40.080 ;
        RECT 1041.050 39.880 1073.570 40.020 ;
        RECT 1041.050 39.820 1041.370 39.880 ;
        RECT 1073.250 39.820 1073.570 39.880 ;
      LAYER via ;
        RECT 1041.080 39.820 1041.340 40.080 ;
        RECT 1073.280 39.820 1073.540 40.080 ;
      LAYER met2 ;
        RECT 1039.650 216.650 1039.930 220.000 ;
        RECT 1039.650 216.510 1041.280 216.650 ;
        RECT 1039.650 216.000 1039.930 216.510 ;
        RECT 1041.140 40.110 1041.280 216.510 ;
        RECT 1041.080 39.790 1041.340 40.110 ;
        RECT 1073.280 39.790 1073.540 40.110 ;
        RECT 1073.340 2.400 1073.480 39.790 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1090.730 43.760 1091.050 43.820 ;
        RECT 1186.870 43.760 1187.190 43.820 ;
        RECT 1090.730 43.620 1187.190 43.760 ;
        RECT 1090.730 43.560 1091.050 43.620 ;
        RECT 1186.870 43.560 1187.190 43.620 ;
      LAYER via ;
        RECT 1090.760 43.560 1091.020 43.820 ;
        RECT 1186.900 43.560 1187.160 43.820 ;
      LAYER met2 ;
        RECT 1187.770 216.650 1188.050 220.000 ;
        RECT 1186.960 216.510 1188.050 216.650 ;
        RECT 1186.960 43.850 1187.100 216.510 ;
        RECT 1187.770 216.000 1188.050 216.510 ;
        RECT 1090.760 43.530 1091.020 43.850 ;
        RECT 1186.900 43.530 1187.160 43.850 ;
        RECT 1090.820 2.400 1090.960 43.530 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 305.510 39.000 305.830 39.060 ;
        RECT 1108.670 39.000 1108.990 39.060 ;
        RECT 305.510 38.860 1108.990 39.000 ;
        RECT 305.510 38.800 305.830 38.860 ;
        RECT 1108.670 38.800 1108.990 38.860 ;
      LAYER via ;
        RECT 305.540 38.800 305.800 39.060 ;
        RECT 1108.700 38.800 1108.960 39.060 ;
      LAYER met2 ;
        RECT 305.530 818.875 305.810 819.245 ;
        RECT 305.600 39.090 305.740 818.875 ;
        RECT 305.540 38.770 305.800 39.090 ;
        RECT 1108.700 38.770 1108.960 39.090 ;
        RECT 1108.760 2.400 1108.900 38.770 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
      LAYER via2 ;
        RECT 305.530 818.920 305.810 819.200 ;
      LAYER met3 ;
        RECT 305.505 819.210 305.835 819.225 ;
        RECT 305.505 819.120 310.500 819.210 ;
        RECT 305.505 818.910 314.000 819.120 ;
        RECT 305.505 818.895 305.835 818.910 ;
        RECT 310.000 818.520 314.000 818.910 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 903.510 46.140 903.830 46.200 ;
        RECT 1126.610 46.140 1126.930 46.200 ;
        RECT 903.510 46.000 1126.930 46.140 ;
        RECT 903.510 45.940 903.830 46.000 ;
        RECT 1126.610 45.940 1126.930 46.000 ;
      LAYER via ;
        RECT 903.540 45.940 903.800 46.200 ;
        RECT 1126.640 45.940 1126.900 46.200 ;
      LAYER met2 ;
        RECT 900.730 216.650 901.010 220.000 ;
        RECT 900.730 216.510 903.740 216.650 ;
        RECT 900.730 216.000 901.010 216.510 ;
        RECT 903.600 46.230 903.740 216.510 ;
        RECT 903.540 45.910 903.800 46.230 ;
        RECT 1126.640 45.910 1126.900 46.230 ;
        RECT 1126.700 2.400 1126.840 45.910 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.410 44.780 634.730 44.840 ;
        RECT 1144.550 44.780 1144.870 44.840 ;
        RECT 634.410 44.640 1144.870 44.780 ;
        RECT 634.410 44.580 634.730 44.640 ;
        RECT 1144.550 44.580 1144.870 44.640 ;
      LAYER via ;
        RECT 634.440 44.580 634.700 44.840 ;
        RECT 1144.580 44.580 1144.840 44.840 ;
      LAYER met2 ;
        RECT 633.930 216.650 634.210 220.000 ;
        RECT 633.930 216.510 634.640 216.650 ;
        RECT 633.930 216.000 634.210 216.510 ;
        RECT 634.500 44.870 634.640 216.510 ;
        RECT 634.440 44.550 634.700 44.870 ;
        RECT 1144.580 44.550 1144.840 44.870 ;
        RECT 1144.640 2.400 1144.780 44.550 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 869.085 1314.865 869.255 1321.495 ;
      LAYER mcon ;
        RECT 869.085 1321.325 869.255 1321.495 ;
      LAYER met1 ;
        RECT 869.010 1321.480 869.330 1321.540 ;
        RECT 868.815 1321.340 869.330 1321.480 ;
        RECT 869.010 1321.280 869.330 1321.340 ;
        RECT 869.025 1315.020 869.315 1315.065 ;
        RECT 1405.370 1315.020 1405.690 1315.080 ;
        RECT 869.025 1314.880 1405.690 1315.020 ;
        RECT 869.025 1314.835 869.315 1314.880 ;
        RECT 1405.370 1314.820 1405.690 1314.880 ;
        RECT 1405.370 484.200 1405.690 484.460 ;
        RECT 1405.460 483.440 1405.600 484.200 ;
        RECT 1405.370 483.180 1405.690 483.440 ;
      LAYER via ;
        RECT 869.040 1321.280 869.300 1321.540 ;
        RECT 1405.400 1314.820 1405.660 1315.080 ;
        RECT 1405.400 484.200 1405.660 484.460 ;
        RECT 1405.400 483.180 1405.660 483.440 ;
      LAYER met2 ;
        RECT 868.530 1321.650 868.810 1325.025 ;
        RECT 868.530 1321.570 869.240 1321.650 ;
        RECT 868.530 1321.510 869.300 1321.570 ;
        RECT 868.530 1321.025 868.810 1321.510 ;
        RECT 869.040 1321.250 869.300 1321.510 ;
        RECT 1405.400 1314.790 1405.660 1315.110 ;
        RECT 1405.460 484.490 1405.600 1314.790 ;
        RECT 1405.400 484.170 1405.660 484.490 ;
        RECT 1405.400 483.150 1405.660 483.470 ;
        RECT 1405.460 304.485 1405.600 483.150 ;
        RECT 1405.390 304.115 1405.670 304.485 ;
        RECT 1162.510 17.835 1162.790 18.205 ;
        RECT 1162.580 2.400 1162.720 17.835 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
      LAYER via2 ;
        RECT 1405.390 304.160 1405.670 304.440 ;
        RECT 1162.510 17.880 1162.790 18.160 ;
      LAYER met3 ;
        RECT 1405.365 304.450 1405.695 304.465 ;
        RECT 1406.950 304.450 1407.330 304.460 ;
        RECT 1405.365 304.150 1407.330 304.450 ;
        RECT 1405.365 304.135 1405.695 304.150 ;
        RECT 1406.950 304.140 1407.330 304.150 ;
        RECT 1162.485 18.170 1162.815 18.185 ;
        RECT 1398.670 18.170 1399.050 18.180 ;
        RECT 1162.485 17.870 1399.050 18.170 ;
        RECT 1162.485 17.855 1162.815 17.870 ;
        RECT 1398.670 17.860 1399.050 17.870 ;
      LAYER via3 ;
        RECT 1406.980 304.140 1407.300 304.460 ;
        RECT 1398.700 17.860 1399.020 18.180 ;
      LAYER met4 ;
        RECT 1398.270 303.710 1399.450 304.890 ;
        RECT 1406.550 303.710 1407.730 304.890 ;
        RECT 1398.710 18.185 1399.010 303.710 ;
        RECT 1398.695 17.855 1399.025 18.185 ;
      LAYER met5 ;
        RECT 1398.060 303.500 1407.940 305.100 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 680.410 17.240 680.730 17.300 ;
        RECT 682.710 17.240 683.030 17.300 ;
        RECT 680.410 17.100 683.030 17.240 ;
        RECT 680.410 17.040 680.730 17.100 ;
        RECT 682.710 17.040 683.030 17.100 ;
      LAYER via ;
        RECT 680.440 17.040 680.700 17.300 ;
        RECT 682.740 17.040 683.000 17.300 ;
      LAYER met2 ;
        RECT 1230.130 1347.915 1230.410 1348.285 ;
        RECT 1230.200 1325.025 1230.340 1347.915 ;
        RECT 1230.090 1321.025 1230.370 1325.025 ;
        RECT 682.730 195.995 683.010 196.365 ;
        RECT 682.800 17.330 682.940 195.995 ;
        RECT 680.440 17.010 680.700 17.330 ;
        RECT 682.740 17.010 683.000 17.330 ;
        RECT 680.500 2.400 680.640 17.010 ;
        RECT 680.290 -4.800 680.850 2.400 ;
      LAYER via2 ;
        RECT 1230.130 1347.960 1230.410 1348.240 ;
        RECT 682.730 196.040 683.010 196.320 ;
      LAYER met3 ;
        RECT 1230.105 1348.250 1230.435 1348.265 ;
        RECT 1402.350 1348.250 1402.730 1348.260 ;
        RECT 1230.105 1347.950 1402.730 1348.250 ;
        RECT 1230.105 1347.935 1230.435 1347.950 ;
        RECT 1402.350 1347.940 1402.730 1347.950 ;
        RECT 682.705 196.330 683.035 196.345 ;
        RECT 1402.350 196.330 1402.730 196.340 ;
        RECT 682.705 196.030 1402.730 196.330 ;
        RECT 682.705 196.015 683.035 196.030 ;
        RECT 1402.350 196.020 1402.730 196.030 ;
      LAYER via3 ;
        RECT 1402.380 1347.940 1402.700 1348.260 ;
        RECT 1402.380 196.020 1402.700 196.340 ;
      LAYER met4 ;
        RECT 1402.375 1347.935 1402.705 1348.265 ;
        RECT 1402.390 196.345 1402.690 1347.935 ;
        RECT 1402.375 196.015 1402.705 196.345 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 305.970 128.080 306.290 128.140 ;
        RECT 1179.970 128.080 1180.290 128.140 ;
        RECT 305.970 127.940 1180.290 128.080 ;
        RECT 305.970 127.880 306.290 127.940 ;
        RECT 1179.970 127.880 1180.290 127.940 ;
      LAYER via ;
        RECT 306.000 127.880 306.260 128.140 ;
        RECT 1180.000 127.880 1180.260 128.140 ;
      LAYER met2 ;
        RECT 305.990 473.435 306.270 473.805 ;
        RECT 306.060 128.170 306.200 473.435 ;
        RECT 306.000 127.850 306.260 128.170 ;
        RECT 1180.000 127.850 1180.260 128.170 ;
        RECT 1180.060 2.400 1180.200 127.850 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
      LAYER via2 ;
        RECT 305.990 473.480 306.270 473.760 ;
      LAYER met3 ;
        RECT 310.000 475.800 314.000 476.400 ;
        RECT 305.965 473.770 306.295 473.785 ;
        RECT 310.350 473.770 310.650 475.800 ;
        RECT 305.965 473.470 310.650 473.770 ;
        RECT 305.965 473.455 306.295 473.470 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1200.210 73.000 1200.530 73.060 ;
        RECT 1406.290 73.000 1406.610 73.060 ;
        RECT 1200.210 72.860 1406.610 73.000 ;
        RECT 1200.210 72.800 1200.530 72.860 ;
        RECT 1406.290 72.800 1406.610 72.860 ;
        RECT 1197.910 20.640 1198.230 20.700 ;
        RECT 1200.210 20.640 1200.530 20.700 ;
        RECT 1197.910 20.500 1200.530 20.640 ;
        RECT 1197.910 20.440 1198.230 20.500 ;
        RECT 1200.210 20.440 1200.530 20.500 ;
      LAYER via ;
        RECT 1200.240 72.800 1200.500 73.060 ;
        RECT 1406.320 72.800 1406.580 73.060 ;
        RECT 1197.940 20.440 1198.200 20.700 ;
        RECT 1200.240 20.440 1200.500 20.700 ;
      LAYER met2 ;
        RECT 1406.310 692.395 1406.590 692.765 ;
        RECT 1406.380 73.090 1406.520 692.395 ;
        RECT 1200.240 72.770 1200.500 73.090 ;
        RECT 1406.320 72.770 1406.580 73.090 ;
        RECT 1200.300 20.730 1200.440 72.770 ;
        RECT 1197.940 20.410 1198.200 20.730 ;
        RECT 1200.240 20.410 1200.500 20.730 ;
        RECT 1198.000 2.400 1198.140 20.410 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
      LAYER via2 ;
        RECT 1406.310 692.440 1406.590 692.720 ;
      LAYER met3 ;
        RECT 1404.305 694.760 1408.305 695.360 ;
        RECT 1406.070 692.745 1406.370 694.760 ;
        RECT 1406.070 692.430 1406.615 692.745 ;
        RECT 1406.285 692.415 1406.615 692.430 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 813.810 47.840 814.130 47.900 ;
        RECT 1215.850 47.840 1216.170 47.900 ;
        RECT 813.810 47.700 1216.170 47.840 ;
        RECT 813.810 47.640 814.130 47.700 ;
        RECT 1215.850 47.640 1216.170 47.700 ;
      LAYER via ;
        RECT 813.840 47.640 814.100 47.900 ;
        RECT 1215.880 47.640 1216.140 47.900 ;
      LAYER met2 ;
        RECT 811.490 216.650 811.770 220.000 ;
        RECT 811.490 216.510 814.040 216.650 ;
        RECT 811.490 216.000 811.770 216.510 ;
        RECT 813.900 47.930 814.040 216.510 ;
        RECT 813.840 47.610 814.100 47.930 ;
        RECT 1215.880 47.610 1216.140 47.930 ;
        RECT 1215.940 2.400 1216.080 47.610 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 293.550 134.880 293.870 134.940 ;
        RECT 1228.730 134.880 1229.050 134.940 ;
        RECT 293.550 134.740 1229.050 134.880 ;
        RECT 293.550 134.680 293.870 134.740 ;
        RECT 1228.730 134.680 1229.050 134.740 ;
      LAYER via ;
        RECT 293.580 134.680 293.840 134.940 ;
        RECT 1228.760 134.680 1229.020 134.940 ;
      LAYER met2 ;
        RECT 293.570 731.835 293.850 732.205 ;
        RECT 293.640 134.970 293.780 731.835 ;
        RECT 293.580 134.650 293.840 134.970 ;
        RECT 1228.760 134.650 1229.020 134.970 ;
        RECT 1228.820 16.730 1228.960 134.650 ;
        RECT 1228.820 16.590 1234.020 16.730 ;
        RECT 1233.880 2.400 1234.020 16.590 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
      LAYER via2 ;
        RECT 293.570 731.880 293.850 732.160 ;
      LAYER met3 ;
        RECT 293.545 732.170 293.875 732.185 ;
        RECT 293.545 732.080 310.500 732.170 ;
        RECT 293.545 731.870 314.000 732.080 ;
        RECT 293.545 731.855 293.875 731.870 ;
        RECT 310.000 731.480 314.000 731.870 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 848.310 48.180 848.630 48.240 ;
        RECT 1251.730 48.180 1252.050 48.240 ;
        RECT 848.310 48.040 1252.050 48.180 ;
        RECT 848.310 47.980 848.630 48.040 ;
        RECT 1251.730 47.980 1252.050 48.040 ;
      LAYER via ;
        RECT 848.340 47.980 848.600 48.240 ;
        RECT 1251.760 47.980 1252.020 48.240 ;
      LAYER met2 ;
        RECT 846.450 216.650 846.730 220.000 ;
        RECT 846.450 216.510 848.540 216.650 ;
        RECT 846.450 216.000 846.730 216.510 ;
        RECT 848.400 48.270 848.540 216.510 ;
        RECT 848.340 47.950 848.600 48.270 ;
        RECT 1251.760 47.950 1252.020 48.270 ;
        RECT 1251.820 2.400 1251.960 47.950 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 294.010 176.700 294.330 176.760 ;
        RECT 1262.770 176.700 1263.090 176.760 ;
        RECT 294.010 176.560 1263.090 176.700 ;
        RECT 294.010 176.500 294.330 176.560 ;
        RECT 1262.770 176.500 1263.090 176.560 ;
        RECT 1262.770 16.900 1263.090 16.960 ;
        RECT 1269.210 16.900 1269.530 16.960 ;
        RECT 1262.770 16.760 1269.530 16.900 ;
        RECT 1262.770 16.700 1263.090 16.760 ;
        RECT 1269.210 16.700 1269.530 16.760 ;
      LAYER via ;
        RECT 294.040 176.500 294.300 176.760 ;
        RECT 1262.800 176.500 1263.060 176.760 ;
        RECT 1262.800 16.700 1263.060 16.960 ;
        RECT 1269.240 16.700 1269.500 16.960 ;
      LAYER met2 ;
        RECT 294.030 870.555 294.310 870.925 ;
        RECT 294.100 176.790 294.240 870.555 ;
        RECT 294.040 176.470 294.300 176.790 ;
        RECT 1262.800 176.470 1263.060 176.790 ;
        RECT 1262.860 16.990 1263.000 176.470 ;
        RECT 1262.800 16.670 1263.060 16.990 ;
        RECT 1269.240 16.670 1269.500 16.990 ;
        RECT 1269.300 2.400 1269.440 16.670 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
      LAYER via2 ;
        RECT 294.030 870.600 294.310 870.880 ;
      LAYER met3 ;
        RECT 294.005 870.890 294.335 870.905 ;
        RECT 294.005 870.800 310.500 870.890 ;
        RECT 294.005 870.590 314.000 870.800 ;
        RECT 294.005 870.575 294.335 870.590 ;
        RECT 310.000 870.200 314.000 870.590 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 893.390 1341.880 893.710 1341.940 ;
        RECT 1443.090 1341.880 1443.410 1341.940 ;
        RECT 893.390 1341.740 1443.410 1341.880 ;
        RECT 893.390 1341.680 893.710 1341.740 ;
        RECT 1443.090 1341.680 1443.410 1341.740 ;
        RECT 1287.150 48.180 1287.470 48.240 ;
        RECT 1443.090 48.180 1443.410 48.240 ;
        RECT 1287.150 48.040 1443.410 48.180 ;
        RECT 1287.150 47.980 1287.470 48.040 ;
        RECT 1443.090 47.980 1443.410 48.040 ;
      LAYER via ;
        RECT 893.420 1341.680 893.680 1341.940 ;
        RECT 1443.120 1341.680 1443.380 1341.940 ;
        RECT 1287.180 47.980 1287.440 48.240 ;
        RECT 1443.120 47.980 1443.380 48.240 ;
      LAYER met2 ;
        RECT 893.420 1341.650 893.680 1341.970 ;
        RECT 1443.120 1341.650 1443.380 1341.970 ;
        RECT 893.480 1325.025 893.620 1341.650 ;
        RECT 893.370 1321.025 893.650 1325.025 ;
        RECT 1443.180 48.270 1443.320 1341.650 ;
        RECT 1287.180 47.950 1287.440 48.270 ;
        RECT 1443.120 47.950 1443.380 48.270 ;
        RECT 1287.240 2.400 1287.380 47.950 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1338.670 1332.360 1338.990 1332.420 ;
        RECT 1443.550 1332.360 1443.870 1332.420 ;
        RECT 1338.670 1332.220 1443.870 1332.360 ;
        RECT 1338.670 1332.160 1338.990 1332.220 ;
        RECT 1443.550 1332.160 1443.870 1332.220 ;
        RECT 1310.610 209.680 1310.930 209.740 ;
        RECT 1443.550 209.680 1443.870 209.740 ;
        RECT 1310.610 209.540 1443.870 209.680 ;
        RECT 1310.610 209.480 1310.930 209.540 ;
        RECT 1443.550 209.480 1443.870 209.540 ;
        RECT 1305.090 16.900 1305.410 16.960 ;
        RECT 1310.610 16.900 1310.930 16.960 ;
        RECT 1305.090 16.760 1310.930 16.900 ;
        RECT 1305.090 16.700 1305.410 16.760 ;
        RECT 1310.610 16.700 1310.930 16.760 ;
      LAYER via ;
        RECT 1338.700 1332.160 1338.960 1332.420 ;
        RECT 1443.580 1332.160 1443.840 1332.420 ;
        RECT 1310.640 209.480 1310.900 209.740 ;
        RECT 1443.580 209.480 1443.840 209.740 ;
        RECT 1305.120 16.700 1305.380 16.960 ;
        RECT 1310.640 16.700 1310.900 16.960 ;
      LAYER met2 ;
        RECT 1338.700 1332.130 1338.960 1332.450 ;
        RECT 1443.580 1332.130 1443.840 1332.450 ;
        RECT 1338.760 1325.025 1338.900 1332.130 ;
        RECT 1338.650 1321.025 1338.930 1325.025 ;
        RECT 1443.640 209.770 1443.780 1332.130 ;
        RECT 1310.640 209.450 1310.900 209.770 ;
        RECT 1443.580 209.450 1443.840 209.770 ;
        RECT 1310.700 16.990 1310.840 209.450 ;
        RECT 1305.120 16.670 1305.380 16.990 ;
        RECT 1310.640 16.670 1310.900 16.990 ;
        RECT 1305.180 2.400 1305.320 16.670 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 938.470 1349.020 938.790 1349.080 ;
        RECT 1449.070 1349.020 1449.390 1349.080 ;
        RECT 938.470 1348.880 1449.390 1349.020 ;
        RECT 938.470 1348.820 938.790 1348.880 ;
        RECT 1449.070 1348.820 1449.390 1348.880 ;
        RECT 1323.030 44.440 1323.350 44.500 ;
        RECT 1449.070 44.440 1449.390 44.500 ;
        RECT 1323.030 44.300 1449.390 44.440 ;
        RECT 1323.030 44.240 1323.350 44.300 ;
        RECT 1449.070 44.240 1449.390 44.300 ;
      LAYER via ;
        RECT 938.500 1348.820 938.760 1349.080 ;
        RECT 1449.100 1348.820 1449.360 1349.080 ;
        RECT 1323.060 44.240 1323.320 44.500 ;
        RECT 1449.100 44.240 1449.360 44.500 ;
      LAYER met2 ;
        RECT 938.500 1348.790 938.760 1349.110 ;
        RECT 1449.100 1348.790 1449.360 1349.110 ;
        RECT 938.560 1325.025 938.700 1348.790 ;
        RECT 938.450 1321.025 938.730 1325.025 ;
        RECT 1449.160 44.530 1449.300 1348.790 ;
        RECT 1323.060 44.210 1323.320 44.530 ;
        RECT 1449.100 44.210 1449.360 44.530 ;
        RECT 1323.120 2.400 1323.260 44.210 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1403.990 859.760 1404.310 859.820 ;
        RECT 1405.830 859.760 1406.150 859.820 ;
        RECT 1403.990 859.620 1406.150 859.760 ;
        RECT 1403.990 859.560 1404.310 859.620 ;
        RECT 1405.830 859.560 1406.150 859.620 ;
        RECT 1403.990 810.800 1404.310 810.860 ;
        RECT 1406.290 810.800 1406.610 810.860 ;
        RECT 1403.990 810.660 1406.610 810.800 ;
        RECT 1403.990 810.600 1404.310 810.660 ;
        RECT 1406.290 810.600 1406.610 810.660 ;
        RECT 1403.990 762.180 1404.310 762.240 ;
        RECT 1406.290 762.180 1406.610 762.240 ;
        RECT 1403.990 762.040 1406.610 762.180 ;
        RECT 1403.990 761.980 1404.310 762.040 ;
        RECT 1406.290 761.980 1406.610 762.040 ;
        RECT 1403.990 627.540 1404.310 627.600 ;
        RECT 1406.750 627.540 1407.070 627.600 ;
        RECT 1403.990 627.400 1407.070 627.540 ;
        RECT 1403.990 627.340 1404.310 627.400 ;
        RECT 1406.750 627.340 1407.070 627.400 ;
        RECT 1403.990 561.920 1404.310 561.980 ;
        RECT 1406.750 561.920 1407.070 561.980 ;
        RECT 1403.990 561.780 1407.070 561.920 ;
        RECT 1403.990 561.720 1404.310 561.780 ;
        RECT 1406.750 561.720 1407.070 561.780 ;
        RECT 1403.990 532.680 1404.310 532.740 ;
        RECT 1406.750 532.680 1407.070 532.740 ;
        RECT 1403.990 532.540 1407.070 532.680 ;
        RECT 1403.990 532.480 1404.310 532.540 ;
        RECT 1406.750 532.480 1407.070 532.540 ;
        RECT 1403.990 472.500 1404.310 472.560 ;
        RECT 1406.750 472.500 1407.070 472.560 ;
        RECT 1403.990 472.360 1407.070 472.500 ;
        RECT 1403.990 472.300 1404.310 472.360 ;
        RECT 1406.750 472.300 1407.070 472.360 ;
        RECT 1403.990 425.240 1404.310 425.300 ;
        RECT 1407.210 425.240 1407.530 425.300 ;
        RECT 1403.990 425.100 1407.530 425.240 ;
        RECT 1403.990 425.040 1404.310 425.100 ;
        RECT 1407.210 425.040 1407.530 425.100 ;
        RECT 1403.990 375.940 1404.310 376.000 ;
        RECT 1407.210 375.940 1407.530 376.000 ;
        RECT 1403.990 375.800 1407.530 375.940 ;
        RECT 1403.990 375.740 1404.310 375.800 ;
        RECT 1407.210 375.740 1407.530 375.800 ;
        RECT 1403.990 337.180 1404.310 337.240 ;
        RECT 1407.210 337.180 1407.530 337.240 ;
        RECT 1403.990 337.040 1407.530 337.180 ;
        RECT 1403.990 336.980 1404.310 337.040 ;
        RECT 1407.210 336.980 1407.530 337.040 ;
        RECT 1407.210 255.580 1407.530 255.640 ;
        RECT 1404.080 255.440 1407.530 255.580 ;
        RECT 1404.080 255.300 1404.220 255.440 ;
        RECT 1407.210 255.380 1407.530 255.440 ;
        RECT 1403.990 255.040 1404.310 255.300 ;
        RECT 1403.990 241.300 1404.310 241.360 ;
        RECT 1406.750 241.300 1407.070 241.360 ;
        RECT 1403.990 241.160 1407.070 241.300 ;
        RECT 1403.990 241.100 1404.310 241.160 ;
        RECT 1406.750 241.100 1407.070 241.160 ;
        RECT 1404.450 182.480 1404.770 182.540 ;
        RECT 1406.750 182.480 1407.070 182.540 ;
        RECT 1404.450 182.340 1407.070 182.480 ;
        RECT 1404.450 182.280 1404.770 182.340 ;
        RECT 1406.750 182.280 1407.070 182.340 ;
        RECT 1345.110 162.420 1345.430 162.480 ;
        RECT 1404.450 162.420 1404.770 162.480 ;
        RECT 1345.110 162.280 1404.770 162.420 ;
        RECT 1345.110 162.220 1345.430 162.280 ;
        RECT 1404.450 162.220 1404.770 162.280 ;
        RECT 1340.510 16.220 1340.830 16.280 ;
        RECT 1345.110 16.220 1345.430 16.280 ;
        RECT 1340.510 16.080 1345.430 16.220 ;
        RECT 1340.510 16.020 1340.830 16.080 ;
        RECT 1345.110 16.020 1345.430 16.080 ;
      LAYER via ;
        RECT 1404.020 859.560 1404.280 859.820 ;
        RECT 1405.860 859.560 1406.120 859.820 ;
        RECT 1404.020 810.600 1404.280 810.860 ;
        RECT 1406.320 810.600 1406.580 810.860 ;
        RECT 1404.020 761.980 1404.280 762.240 ;
        RECT 1406.320 761.980 1406.580 762.240 ;
        RECT 1404.020 627.340 1404.280 627.600 ;
        RECT 1406.780 627.340 1407.040 627.600 ;
        RECT 1404.020 561.720 1404.280 561.980 ;
        RECT 1406.780 561.720 1407.040 561.980 ;
        RECT 1404.020 532.480 1404.280 532.740 ;
        RECT 1406.780 532.480 1407.040 532.740 ;
        RECT 1404.020 472.300 1404.280 472.560 ;
        RECT 1406.780 472.300 1407.040 472.560 ;
        RECT 1404.020 425.040 1404.280 425.300 ;
        RECT 1407.240 425.040 1407.500 425.300 ;
        RECT 1404.020 375.740 1404.280 376.000 ;
        RECT 1407.240 375.740 1407.500 376.000 ;
        RECT 1404.020 336.980 1404.280 337.240 ;
        RECT 1407.240 336.980 1407.500 337.240 ;
        RECT 1407.240 255.380 1407.500 255.640 ;
        RECT 1404.020 255.040 1404.280 255.300 ;
        RECT 1404.020 241.100 1404.280 241.360 ;
        RECT 1406.780 241.100 1407.040 241.360 ;
        RECT 1404.480 182.280 1404.740 182.540 ;
        RECT 1406.780 182.280 1407.040 182.540 ;
        RECT 1345.140 162.220 1345.400 162.480 ;
        RECT 1404.480 162.220 1404.740 162.480 ;
        RECT 1340.540 16.020 1340.800 16.280 ;
        RECT 1345.140 16.020 1345.400 16.280 ;
      LAYER met2 ;
        RECT 1405.850 948.075 1406.130 948.445 ;
        RECT 1405.920 859.850 1406.060 948.075 ;
        RECT 1404.020 859.530 1404.280 859.850 ;
        RECT 1405.860 859.530 1406.120 859.850 ;
        RECT 1404.080 810.890 1404.220 859.530 ;
        RECT 1404.020 810.570 1404.280 810.890 ;
        RECT 1406.320 810.570 1406.580 810.890 ;
        RECT 1406.380 762.270 1406.520 810.570 ;
        RECT 1404.020 761.950 1404.280 762.270 ;
        RECT 1406.320 761.950 1406.580 762.270 ;
        RECT 1404.080 627.630 1404.220 761.950 ;
        RECT 1404.020 627.310 1404.280 627.630 ;
        RECT 1406.780 627.310 1407.040 627.630 ;
        RECT 1406.840 562.010 1406.980 627.310 ;
        RECT 1404.020 561.690 1404.280 562.010 ;
        RECT 1406.780 561.690 1407.040 562.010 ;
        RECT 1404.080 532.770 1404.220 561.690 ;
        RECT 1404.020 532.450 1404.280 532.770 ;
        RECT 1406.780 532.450 1407.040 532.770 ;
        RECT 1406.840 472.590 1406.980 532.450 ;
        RECT 1404.020 472.270 1404.280 472.590 ;
        RECT 1406.780 472.270 1407.040 472.590 ;
        RECT 1404.080 425.330 1404.220 472.270 ;
        RECT 1404.020 425.010 1404.280 425.330 ;
        RECT 1407.240 425.010 1407.500 425.330 ;
        RECT 1407.300 376.030 1407.440 425.010 ;
        RECT 1404.020 375.710 1404.280 376.030 ;
        RECT 1407.240 375.710 1407.500 376.030 ;
        RECT 1404.080 337.270 1404.220 375.710 ;
        RECT 1404.020 336.950 1404.280 337.270 ;
        RECT 1407.240 336.950 1407.500 337.270 ;
        RECT 1407.300 255.670 1407.440 336.950 ;
        RECT 1407.240 255.350 1407.500 255.670 ;
        RECT 1404.020 255.010 1404.280 255.330 ;
        RECT 1404.080 241.390 1404.220 255.010 ;
        RECT 1404.020 241.070 1404.280 241.390 ;
        RECT 1406.780 241.070 1407.040 241.390 ;
        RECT 1406.840 182.570 1406.980 241.070 ;
        RECT 1404.480 182.250 1404.740 182.570 ;
        RECT 1406.780 182.250 1407.040 182.570 ;
        RECT 1404.540 162.510 1404.680 182.250 ;
        RECT 1345.140 162.190 1345.400 162.510 ;
        RECT 1404.480 162.190 1404.740 162.510 ;
        RECT 1345.200 16.310 1345.340 162.190 ;
        RECT 1340.540 15.990 1340.800 16.310 ;
        RECT 1345.140 15.990 1345.400 16.310 ;
        RECT 1340.600 2.400 1340.740 15.990 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
      LAYER via2 ;
        RECT 1405.850 948.120 1406.130 948.400 ;
      LAYER met3 ;
        RECT 1404.305 950.440 1408.305 951.040 ;
        RECT 1406.070 948.425 1406.370 950.440 ;
        RECT 1405.825 948.110 1406.370 948.425 ;
        RECT 1405.825 948.095 1406.155 948.110 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 15.795 698.650 16.165 ;
        RECT 698.440 2.400 698.580 15.795 ;
        RECT 698.230 -4.800 698.790 2.400 ;
      LAYER via2 ;
        RECT 698.370 15.840 698.650 16.120 ;
      LAYER met3 ;
        RECT 300.190 548.570 300.570 548.580 ;
        RECT 300.190 548.480 310.500 548.570 ;
        RECT 300.190 548.270 314.000 548.480 ;
        RECT 300.190 548.260 300.570 548.270 ;
        RECT 310.000 547.880 314.000 548.270 ;
        RECT 318.590 16.130 318.970 16.140 ;
        RECT 698.345 16.130 698.675 16.145 ;
        RECT 318.590 15.830 698.675 16.130 ;
        RECT 318.590 15.820 318.970 15.830 ;
        RECT 698.345 15.815 698.675 15.830 ;
      LAYER via3 ;
        RECT 300.220 548.260 300.540 548.580 ;
        RECT 318.620 15.820 318.940 16.140 ;
      LAYER met4 ;
        RECT 300.215 548.255 300.545 548.585 ;
        RECT 300.230 345.690 300.530 548.255 ;
        RECT 299.790 344.510 300.970 345.690 ;
        RECT 318.190 344.510 319.370 345.690 ;
        RECT 318.630 260.250 318.930 344.510 ;
        RECT 317.710 259.950 318.930 260.250 ;
        RECT 317.710 246.650 318.010 259.950 ;
        RECT 317.710 246.350 318.930 246.650 ;
        RECT 318.630 16.145 318.930 246.350 ;
        RECT 318.615 15.815 318.945 16.145 ;
      LAYER met5 ;
        RECT 299.580 344.300 319.580 345.900 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1338.210 25.400 1338.530 25.460 ;
        RECT 1358.450 25.400 1358.770 25.460 ;
        RECT 1338.210 25.260 1358.770 25.400 ;
        RECT 1338.210 25.200 1338.530 25.260 ;
        RECT 1358.450 25.200 1358.770 25.260 ;
      LAYER via ;
        RECT 1338.240 25.200 1338.500 25.460 ;
        RECT 1358.480 25.200 1358.740 25.460 ;
      LAYER met2 ;
        RECT 1335.890 216.650 1336.170 220.000 ;
        RECT 1335.890 216.510 1338.440 216.650 ;
        RECT 1335.890 216.000 1336.170 216.510 ;
        RECT 1338.300 25.490 1338.440 216.510 ;
        RECT 1338.240 25.170 1338.500 25.490 ;
        RECT 1358.480 25.170 1358.740 25.490 ;
        RECT 1358.540 2.400 1358.680 25.170 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 613.710 47.160 614.030 47.220 ;
        RECT 1376.390 47.160 1376.710 47.220 ;
        RECT 613.710 47.020 1376.710 47.160 ;
        RECT 613.710 46.960 614.030 47.020 ;
        RECT 1376.390 46.960 1376.710 47.020 ;
      LAYER via ;
        RECT 613.740 46.960 614.000 47.220 ;
        RECT 1376.420 46.960 1376.680 47.220 ;
      LAYER met2 ;
        RECT 613.690 216.000 613.970 220.000 ;
        RECT 613.800 47.250 613.940 216.000 ;
        RECT 613.740 46.930 614.000 47.250 ;
        RECT 1376.420 46.930 1376.680 47.250 ;
        RECT 1376.480 2.400 1376.620 46.930 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 266.870 1028.400 267.190 1028.460 ;
        RECT 296.770 1028.400 297.090 1028.460 ;
        RECT 266.870 1028.260 297.090 1028.400 ;
        RECT 266.870 1028.200 267.190 1028.260 ;
        RECT 296.770 1028.200 297.090 1028.260 ;
        RECT 266.870 46.480 267.190 46.540 ;
        RECT 1394.330 46.480 1394.650 46.540 ;
        RECT 266.870 46.340 1394.650 46.480 ;
        RECT 266.870 46.280 267.190 46.340 ;
        RECT 1394.330 46.280 1394.650 46.340 ;
      LAYER via ;
        RECT 266.900 1028.200 267.160 1028.460 ;
        RECT 296.800 1028.200 297.060 1028.460 ;
        RECT 266.900 46.280 267.160 46.540 ;
        RECT 1394.360 46.280 1394.620 46.540 ;
      LAYER met2 ;
        RECT 296.790 1031.035 297.070 1031.405 ;
        RECT 296.860 1028.490 297.000 1031.035 ;
        RECT 266.900 1028.170 267.160 1028.490 ;
        RECT 296.800 1028.170 297.060 1028.490 ;
        RECT 266.960 46.570 267.100 1028.170 ;
        RECT 266.900 46.250 267.160 46.570 ;
        RECT 1394.360 46.250 1394.620 46.570 ;
        RECT 1394.420 2.400 1394.560 46.250 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
      LAYER via2 ;
        RECT 296.790 1031.080 297.070 1031.360 ;
      LAYER met3 ;
        RECT 296.765 1031.370 297.095 1031.385 ;
        RECT 296.765 1031.280 310.500 1031.370 ;
        RECT 296.765 1031.070 314.000 1031.280 ;
        RECT 296.765 1031.055 297.095 1031.070 ;
        RECT 310.000 1030.680 314.000 1031.070 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 292.170 614.620 292.490 614.680 ;
        RECT 301.370 614.620 301.690 614.680 ;
        RECT 292.170 614.480 301.690 614.620 ;
        RECT 292.170 614.420 292.490 614.480 ;
        RECT 301.370 614.420 301.690 614.480 ;
        RECT 292.170 183.160 292.490 183.220 ;
        RECT 1407.670 183.160 1407.990 183.220 ;
        RECT 292.170 183.020 1407.990 183.160 ;
        RECT 292.170 182.960 292.490 183.020 ;
        RECT 1407.670 182.960 1407.990 183.020 ;
        RECT 1407.670 20.980 1407.990 21.040 ;
        RECT 1412.270 20.980 1412.590 21.040 ;
        RECT 1407.670 20.840 1412.590 20.980 ;
        RECT 1407.670 20.780 1407.990 20.840 ;
        RECT 1412.270 20.780 1412.590 20.840 ;
      LAYER via ;
        RECT 292.200 614.420 292.460 614.680 ;
        RECT 301.400 614.420 301.660 614.680 ;
        RECT 292.200 182.960 292.460 183.220 ;
        RECT 1407.700 182.960 1407.960 183.220 ;
        RECT 1407.700 20.780 1407.960 21.040 ;
        RECT 1412.300 20.780 1412.560 21.040 ;
      LAYER met2 ;
        RECT 301.390 614.875 301.670 615.245 ;
        RECT 301.460 614.710 301.600 614.875 ;
        RECT 292.200 614.390 292.460 614.710 ;
        RECT 301.400 614.390 301.660 614.710 ;
        RECT 292.260 183.250 292.400 614.390 ;
        RECT 292.200 182.930 292.460 183.250 ;
        RECT 1407.700 182.930 1407.960 183.250 ;
        RECT 1407.760 21.070 1407.900 182.930 ;
        RECT 1407.700 20.750 1407.960 21.070 ;
        RECT 1412.300 20.750 1412.560 21.070 ;
        RECT 1412.360 2.400 1412.500 20.750 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
      LAYER via2 ;
        RECT 301.390 614.920 301.670 615.200 ;
      LAYER met3 ;
        RECT 301.365 615.210 301.695 615.225 ;
        RECT 301.365 615.120 310.500 615.210 ;
        RECT 301.365 614.910 314.000 615.120 ;
        RECT 301.365 614.895 301.695 614.910 ;
        RECT 310.000 614.520 314.000 614.910 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 399.315 311.790 399.685 ;
        RECT 311.580 339.165 311.720 399.315 ;
        RECT 311.510 338.795 311.790 339.165 ;
        RECT 1429.770 189.195 1430.050 189.565 ;
        RECT 1429.840 2.400 1429.980 189.195 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
      LAYER via2 ;
        RECT 311.510 399.360 311.790 399.640 ;
        RECT 311.510 338.840 311.790 339.120 ;
        RECT 1429.770 189.240 1430.050 189.520 ;
      LAYER met3 ;
        RECT 310.000 789.960 314.000 790.560 ;
        RECT 313.110 785.900 313.410 789.960 ;
        RECT 313.070 785.580 313.450 785.900 ;
        RECT 311.230 640.370 311.610 640.380 ;
        RECT 313.070 640.370 313.450 640.380 ;
        RECT 311.230 640.070 313.450 640.370 ;
        RECT 311.230 640.060 311.610 640.070 ;
        RECT 313.070 640.060 313.450 640.070 ;
        RECT 311.230 586.650 311.610 586.660 ;
        RECT 313.070 586.650 313.450 586.660 ;
        RECT 311.230 586.350 313.450 586.650 ;
        RECT 311.230 586.340 311.610 586.350 ;
        RECT 313.070 586.340 313.450 586.350 ;
        RECT 311.485 399.650 311.815 399.665 ;
        RECT 313.070 399.650 313.450 399.660 ;
        RECT 311.485 399.350 313.450 399.650 ;
        RECT 311.485 399.335 311.815 399.350 ;
        RECT 313.070 399.340 313.450 399.350 ;
        RECT 311.485 339.130 311.815 339.145 ;
        RECT 313.070 339.130 313.450 339.140 ;
        RECT 311.485 338.830 313.450 339.130 ;
        RECT 311.485 338.815 311.815 338.830 ;
        RECT 313.070 338.820 313.450 338.830 ;
        RECT 312.150 189.530 312.530 189.540 ;
        RECT 1429.745 189.530 1430.075 189.545 ;
        RECT 312.150 189.230 1430.075 189.530 ;
        RECT 312.150 189.220 312.530 189.230 ;
        RECT 1429.745 189.215 1430.075 189.230 ;
      LAYER via3 ;
        RECT 313.100 785.580 313.420 785.900 ;
        RECT 311.260 640.060 311.580 640.380 ;
        RECT 313.100 640.060 313.420 640.380 ;
        RECT 311.260 586.340 311.580 586.660 ;
        RECT 313.100 586.340 313.420 586.660 ;
        RECT 313.100 399.340 313.420 399.660 ;
        RECT 313.100 338.820 313.420 339.140 ;
        RECT 312.180 189.220 312.500 189.540 ;
      LAYER met4 ;
        RECT 313.095 785.575 313.425 785.905 ;
        RECT 313.110 719.250 313.410 785.575 ;
        RECT 313.110 718.950 315.250 719.250 ;
        RECT 314.950 675.730 315.250 718.950 ;
        RECT 313.110 675.430 315.250 675.730 ;
        RECT 313.110 640.385 313.410 675.430 ;
        RECT 311.255 640.055 311.585 640.385 ;
        RECT 313.095 640.055 313.425 640.385 ;
        RECT 311.270 586.665 311.570 640.055 ;
        RECT 311.255 586.335 311.585 586.665 ;
        RECT 313.095 586.650 313.425 586.665 ;
        RECT 313.095 586.350 316.170 586.650 ;
        RECT 313.095 586.335 313.425 586.350 ;
        RECT 315.870 579.850 316.170 586.350 ;
        RECT 314.030 579.550 316.170 579.850 ;
        RECT 314.030 552.650 314.330 579.550 ;
        RECT 312.190 552.350 314.330 552.650 ;
        RECT 312.190 467.650 312.490 552.350 ;
        RECT 312.190 467.350 316.170 467.650 ;
        RECT 315.870 440.450 316.170 467.350 ;
        RECT 314.030 440.150 316.170 440.450 ;
        RECT 313.095 399.650 313.425 399.665 ;
        RECT 314.030 399.650 314.330 440.150 ;
        RECT 313.095 399.350 314.330 399.650 ;
        RECT 313.095 399.335 313.425 399.350 ;
        RECT 313.095 338.815 313.425 339.145 ;
        RECT 313.110 328.250 313.410 338.815 ;
        RECT 313.110 327.950 314.330 328.250 ;
        RECT 314.030 304.450 314.330 327.950 ;
        RECT 314.030 304.150 316.170 304.450 ;
        RECT 315.870 273.850 316.170 304.150 ;
        RECT 314.030 273.550 316.170 273.850 ;
        RECT 314.030 239.850 314.330 273.550 ;
        RECT 312.190 239.550 314.330 239.850 ;
        RECT 312.190 189.545 312.490 239.550 ;
        RECT 312.175 189.215 312.505 189.545 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1299.110 1336.440 1299.430 1336.500 ;
        RECT 1406.750 1336.440 1407.070 1336.500 ;
        RECT 1299.110 1336.300 1407.070 1336.440 ;
        RECT 1299.110 1336.240 1299.430 1336.300 ;
        RECT 1406.750 1336.240 1407.070 1336.300 ;
        RECT 1406.750 1317.740 1407.070 1317.800 ;
        RECT 1442.170 1317.740 1442.490 1317.800 ;
        RECT 1406.750 1317.600 1442.490 1317.740 ;
        RECT 1406.750 1317.540 1407.070 1317.600 ;
        RECT 1442.170 1317.540 1442.490 1317.600 ;
      LAYER via ;
        RECT 1299.140 1336.240 1299.400 1336.500 ;
        RECT 1406.780 1336.240 1407.040 1336.500 ;
        RECT 1406.780 1317.540 1407.040 1317.800 ;
        RECT 1442.200 1317.540 1442.460 1317.800 ;
      LAYER met2 ;
        RECT 1299.140 1336.210 1299.400 1336.530 ;
        RECT 1406.780 1336.210 1407.040 1336.530 ;
        RECT 1299.200 1325.025 1299.340 1336.210 ;
        RECT 1299.090 1321.025 1299.370 1325.025 ;
        RECT 1406.840 1317.830 1406.980 1336.210 ;
        RECT 1406.780 1317.510 1407.040 1317.830 ;
        RECT 1442.200 1317.510 1442.460 1317.830 ;
        RECT 1442.260 17.410 1442.400 1317.510 ;
        RECT 1442.260 17.270 1447.920 17.410 ;
        RECT 1447.780 2.400 1447.920 17.270 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 911.100 1421.330 911.160 ;
        RECT 1462.870 911.100 1463.190 911.160 ;
        RECT 1421.010 910.960 1463.190 911.100 ;
        RECT 1421.010 910.900 1421.330 910.960 ;
        RECT 1462.870 910.900 1463.190 910.960 ;
      LAYER via ;
        RECT 1421.040 910.900 1421.300 911.160 ;
        RECT 1462.900 910.900 1463.160 911.160 ;
      LAYER met2 ;
        RECT 1421.030 914.075 1421.310 914.445 ;
        RECT 1421.100 911.190 1421.240 914.075 ;
        RECT 1421.040 910.870 1421.300 911.190 ;
        RECT 1462.900 910.870 1463.160 911.190 ;
        RECT 1462.960 16.730 1463.100 910.870 ;
        RECT 1462.960 16.590 1465.860 16.730 ;
        RECT 1465.720 2.400 1465.860 16.590 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
      LAYER via2 ;
        RECT 1421.030 914.120 1421.310 914.400 ;
      LAYER met3 ;
        RECT 1421.005 914.410 1421.335 914.425 ;
        RECT 1408.060 914.320 1421.335 914.410 ;
        RECT 1404.305 914.110 1421.335 914.320 ;
        RECT 1404.305 913.720 1408.305 914.110 ;
        RECT 1421.005 914.095 1421.335 914.110 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.070 1333.040 621.390 1333.100 ;
        RECT 1411.810 1333.040 1412.130 1333.100 ;
        RECT 621.070 1332.900 1412.130 1333.040 ;
        RECT 621.070 1332.840 621.390 1332.900 ;
        RECT 1411.810 1332.840 1412.130 1332.900 ;
        RECT 1411.810 1308.220 1412.130 1308.280 ;
        RECT 1484.030 1308.220 1484.350 1308.280 ;
        RECT 1411.810 1308.080 1484.350 1308.220 ;
        RECT 1411.810 1308.020 1412.130 1308.080 ;
        RECT 1484.030 1308.020 1484.350 1308.080 ;
      LAYER via ;
        RECT 621.100 1332.840 621.360 1333.100 ;
        RECT 1411.840 1332.840 1412.100 1333.100 ;
        RECT 1411.840 1308.020 1412.100 1308.280 ;
        RECT 1484.060 1308.020 1484.320 1308.280 ;
      LAYER met2 ;
        RECT 621.100 1332.810 621.360 1333.130 ;
        RECT 1411.840 1332.810 1412.100 1333.130 ;
        RECT 621.160 1325.025 621.300 1332.810 ;
        RECT 621.050 1321.025 621.330 1325.025 ;
        RECT 1411.900 1308.310 1412.040 1332.810 ;
        RECT 1411.840 1307.990 1412.100 1308.310 ;
        RECT 1484.060 1307.990 1484.320 1308.310 ;
        RECT 1484.120 7.210 1484.260 1307.990 ;
        RECT 1483.660 7.070 1484.260 7.210 ;
        RECT 1483.660 2.400 1483.800 7.070 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 303.670 59.060 303.990 59.120 ;
        RECT 1497.370 59.060 1497.690 59.120 ;
        RECT 303.670 58.920 1497.690 59.060 ;
        RECT 303.670 58.860 303.990 58.920 ;
        RECT 1497.370 58.860 1497.690 58.920 ;
      LAYER via ;
        RECT 303.700 58.860 303.960 59.120 ;
        RECT 1497.400 58.860 1497.660 59.120 ;
      LAYER met2 ;
        RECT 303.690 1264.955 303.970 1265.325 ;
        RECT 303.760 59.150 303.900 1264.955 ;
        RECT 303.700 58.830 303.960 59.150 ;
        RECT 1497.400 58.830 1497.660 59.150 ;
        RECT 1497.460 17.410 1497.600 58.830 ;
        RECT 1497.460 17.270 1501.740 17.410 ;
        RECT 1501.600 2.400 1501.740 17.270 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
      LAYER via2 ;
        RECT 303.690 1265.000 303.970 1265.280 ;
      LAYER met3 ;
        RECT 303.665 1265.290 303.995 1265.305 ;
        RECT 303.665 1265.200 310.500 1265.290 ;
        RECT 303.665 1264.990 314.000 1265.200 ;
        RECT 303.665 1264.975 303.995 1264.990 ;
        RECT 310.000 1264.600 314.000 1264.990 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1222.750 200.500 1223.070 200.560 ;
        RECT 1227.350 200.500 1227.670 200.560 ;
        RECT 1222.750 200.360 1227.670 200.500 ;
        RECT 1222.750 200.300 1223.070 200.360 ;
        RECT 1227.350 200.300 1227.670 200.360 ;
        RECT 1227.350 47.840 1227.670 47.900 ;
        RECT 1518.990 47.840 1519.310 47.900 ;
        RECT 1227.350 47.700 1519.310 47.840 ;
        RECT 1227.350 47.640 1227.670 47.700 ;
        RECT 1518.990 47.640 1519.310 47.700 ;
      LAYER via ;
        RECT 1222.780 200.300 1223.040 200.560 ;
        RECT 1227.380 200.300 1227.640 200.560 ;
        RECT 1227.380 47.640 1227.640 47.900 ;
        RECT 1519.020 47.640 1519.280 47.900 ;
      LAYER met2 ;
        RECT 1222.730 216.000 1223.010 220.000 ;
        RECT 1222.840 200.590 1222.980 216.000 ;
        RECT 1222.780 200.270 1223.040 200.590 ;
        RECT 1227.380 200.270 1227.640 200.590 ;
        RECT 1227.440 47.930 1227.580 200.270 ;
        RECT 1227.380 47.610 1227.640 47.930 ;
        RECT 1519.020 47.610 1519.280 47.930 ;
        RECT 1519.080 2.400 1519.220 47.610 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 716.750 94.080 717.070 94.140 ;
        RECT 1408.130 94.080 1408.450 94.140 ;
        RECT 716.750 93.940 1408.450 94.080 ;
        RECT 716.750 93.880 717.070 93.940 ;
        RECT 1408.130 93.880 1408.450 93.940 ;
      LAYER via ;
        RECT 716.780 93.880 717.040 94.140 ;
        RECT 1408.160 93.880 1408.420 94.140 ;
      LAYER met2 ;
        RECT 1408.150 524.435 1408.430 524.805 ;
        RECT 1408.220 94.170 1408.360 524.435 ;
        RECT 716.780 93.850 717.040 94.170 ;
        RECT 1408.160 93.850 1408.420 94.170 ;
        RECT 716.840 17.410 716.980 93.850 ;
        RECT 716.380 17.270 716.980 17.410 ;
        RECT 716.380 2.400 716.520 17.270 ;
        RECT 716.170 -4.800 716.730 2.400 ;
      LAYER via2 ;
        RECT 1408.150 524.480 1408.430 524.760 ;
      LAYER met3 ;
        RECT 1404.305 526.120 1408.305 526.720 ;
        RECT 1407.910 524.785 1408.210 526.120 ;
        RECT 1407.910 524.470 1408.455 524.785 ;
        RECT 1408.125 524.455 1408.455 524.470 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1284.390 1333.380 1284.710 1333.440 ;
        RECT 1415.490 1333.380 1415.810 1333.440 ;
        RECT 1284.390 1333.240 1415.810 1333.380 ;
        RECT 1284.390 1333.180 1284.710 1333.240 ;
        RECT 1415.490 1333.180 1415.810 1333.240 ;
        RECT 1415.490 1293.940 1415.810 1294.000 ;
        RECT 1531.870 1293.940 1532.190 1294.000 ;
        RECT 1415.490 1293.800 1532.190 1293.940 ;
        RECT 1415.490 1293.740 1415.810 1293.800 ;
        RECT 1531.870 1293.740 1532.190 1293.800 ;
      LAYER via ;
        RECT 1284.420 1333.180 1284.680 1333.440 ;
        RECT 1415.520 1333.180 1415.780 1333.440 ;
        RECT 1415.520 1293.740 1415.780 1294.000 ;
        RECT 1531.900 1293.740 1532.160 1294.000 ;
      LAYER met2 ;
        RECT 1284.420 1333.150 1284.680 1333.470 ;
        RECT 1415.520 1333.150 1415.780 1333.470 ;
        RECT 1284.480 1325.025 1284.620 1333.150 ;
        RECT 1284.370 1321.025 1284.650 1325.025 ;
        RECT 1415.580 1294.030 1415.720 1333.150 ;
        RECT 1415.520 1293.710 1415.780 1294.030 ;
        RECT 1531.900 1293.710 1532.160 1294.030 ;
        RECT 1531.960 17.410 1532.100 1293.710 ;
        RECT 1531.960 17.270 1537.160 17.410 ;
        RECT 1537.020 2.400 1537.160 17.270 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1130.750 1334.400 1131.070 1334.460 ;
        RECT 1438.950 1334.400 1439.270 1334.460 ;
        RECT 1130.750 1334.260 1439.270 1334.400 ;
        RECT 1130.750 1334.200 1131.070 1334.260 ;
        RECT 1438.950 1334.200 1439.270 1334.260 ;
        RECT 1438.950 224.300 1439.270 224.360 ;
        RECT 1552.570 224.300 1552.890 224.360 ;
        RECT 1438.950 224.160 1552.890 224.300 ;
        RECT 1438.950 224.100 1439.270 224.160 ;
        RECT 1552.570 224.100 1552.890 224.160 ;
      LAYER via ;
        RECT 1130.780 1334.200 1131.040 1334.460 ;
        RECT 1438.980 1334.200 1439.240 1334.460 ;
        RECT 1438.980 224.100 1439.240 224.360 ;
        RECT 1552.600 224.100 1552.860 224.360 ;
      LAYER met2 ;
        RECT 1130.780 1334.170 1131.040 1334.490 ;
        RECT 1438.980 1334.170 1439.240 1334.490 ;
        RECT 1130.840 1325.025 1130.980 1334.170 ;
        RECT 1130.730 1321.025 1131.010 1325.025 ;
        RECT 1439.040 224.390 1439.180 1334.170 ;
        RECT 1438.980 224.070 1439.240 224.390 ;
        RECT 1552.600 224.070 1552.860 224.390 ;
        RECT 1552.660 17.410 1552.800 224.070 ;
        RECT 1552.660 17.270 1555.100 17.410 ;
        RECT 1554.960 2.400 1555.100 17.270 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 517.720 1419.490 517.780 ;
        RECT 1566.370 517.720 1566.690 517.780 ;
        RECT 1419.170 517.580 1566.690 517.720 ;
        RECT 1419.170 517.520 1419.490 517.580 ;
        RECT 1566.370 517.520 1566.690 517.580 ;
        RECT 1566.370 16.900 1566.690 16.960 ;
        RECT 1572.810 16.900 1573.130 16.960 ;
        RECT 1566.370 16.760 1573.130 16.900 ;
        RECT 1566.370 16.700 1566.690 16.760 ;
        RECT 1572.810 16.700 1573.130 16.760 ;
      LAYER via ;
        RECT 1419.200 517.520 1419.460 517.780 ;
        RECT 1566.400 517.520 1566.660 517.780 ;
        RECT 1566.400 16.700 1566.660 16.960 ;
        RECT 1572.840 16.700 1573.100 16.960 ;
      LAYER met2 ;
        RECT 1419.190 519.675 1419.470 520.045 ;
        RECT 1419.260 517.810 1419.400 519.675 ;
        RECT 1419.200 517.490 1419.460 517.810 ;
        RECT 1566.400 517.490 1566.660 517.810 ;
        RECT 1566.460 16.990 1566.600 517.490 ;
        RECT 1566.400 16.670 1566.660 16.990 ;
        RECT 1572.840 16.670 1573.100 16.990 ;
        RECT 1572.900 2.400 1573.040 16.670 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
      LAYER via2 ;
        RECT 1419.190 519.720 1419.470 520.000 ;
      LAYER met3 ;
        RECT 1419.165 520.010 1419.495 520.025 ;
        RECT 1408.060 519.920 1419.495 520.010 ;
        RECT 1404.305 519.710 1419.495 519.920 ;
        RECT 1404.305 519.320 1408.305 519.710 ;
        RECT 1419.165 519.695 1419.495 519.710 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 938.010 47.500 938.330 47.560 ;
        RECT 1590.290 47.500 1590.610 47.560 ;
        RECT 938.010 47.360 1590.610 47.500 ;
        RECT 938.010 47.300 938.330 47.360 ;
        RECT 1590.290 47.300 1590.610 47.360 ;
      LAYER via ;
        RECT 938.040 47.300 938.300 47.560 ;
        RECT 1590.320 47.300 1590.580 47.560 ;
      LAYER met2 ;
        RECT 935.690 216.650 935.970 220.000 ;
        RECT 935.690 216.510 938.240 216.650 ;
        RECT 935.690 216.000 935.970 216.510 ;
        RECT 938.100 47.590 938.240 216.510 ;
        RECT 938.040 47.270 938.300 47.590 ;
        RECT 1590.320 47.270 1590.580 47.590 ;
        RECT 1590.380 2.400 1590.520 47.270 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 565.410 46.820 565.730 46.880 ;
        RECT 1608.230 46.820 1608.550 46.880 ;
        RECT 565.410 46.680 1608.550 46.820 ;
        RECT 565.410 46.620 565.730 46.680 ;
        RECT 1608.230 46.620 1608.550 46.680 ;
      LAYER via ;
        RECT 565.440 46.620 565.700 46.880 ;
        RECT 1608.260 46.620 1608.520 46.880 ;
      LAYER met2 ;
        RECT 564.930 216.650 565.210 220.000 ;
        RECT 564.930 216.510 565.640 216.650 ;
        RECT 564.930 216.000 565.210 216.510 ;
        RECT 565.500 46.910 565.640 216.510 ;
        RECT 565.440 46.590 565.700 46.910 ;
        RECT 1608.260 46.590 1608.520 46.910 ;
        RECT 1608.320 2.400 1608.460 46.590 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.130 114.140 304.450 114.200 ;
        RECT 1621.570 114.140 1621.890 114.200 ;
        RECT 304.130 114.000 1621.890 114.140 ;
        RECT 304.130 113.940 304.450 114.000 ;
        RECT 1621.570 113.940 1621.890 114.000 ;
        RECT 1621.570 2.960 1621.890 3.020 ;
        RECT 1626.170 2.960 1626.490 3.020 ;
        RECT 1621.570 2.820 1626.490 2.960 ;
        RECT 1621.570 2.760 1621.890 2.820 ;
        RECT 1626.170 2.760 1626.490 2.820 ;
      LAYER via ;
        RECT 304.160 113.940 304.420 114.200 ;
        RECT 1621.600 113.940 1621.860 114.200 ;
        RECT 1621.600 2.760 1621.860 3.020 ;
        RECT 1626.200 2.760 1626.460 3.020 ;
      LAYER met2 ;
        RECT 304.150 1249.995 304.430 1250.365 ;
        RECT 304.220 114.230 304.360 1249.995 ;
        RECT 304.160 113.910 304.420 114.230 ;
        RECT 1621.600 113.910 1621.860 114.230 ;
        RECT 1621.660 3.050 1621.800 113.910 ;
        RECT 1621.600 2.730 1621.860 3.050 ;
        RECT 1626.200 2.730 1626.460 3.050 ;
        RECT 1626.260 2.400 1626.400 2.730 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
      LAYER via2 ;
        RECT 304.150 1250.040 304.430 1250.320 ;
      LAYER met3 ;
        RECT 304.125 1250.330 304.455 1250.345 ;
        RECT 304.125 1250.240 310.500 1250.330 ;
        RECT 304.125 1250.030 314.000 1250.240 ;
        RECT 304.125 1250.015 304.455 1250.030 ;
        RECT 310.000 1249.640 314.000 1250.030 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 303.210 51.580 303.530 51.640 ;
        RECT 1642.270 51.580 1642.590 51.640 ;
        RECT 303.210 51.440 1642.590 51.580 ;
        RECT 303.210 51.380 303.530 51.440 ;
        RECT 1642.270 51.380 1642.590 51.440 ;
      LAYER via ;
        RECT 303.240 51.380 303.500 51.640 ;
        RECT 1642.300 51.380 1642.560 51.640 ;
      LAYER met2 ;
        RECT 303.230 534.635 303.510 535.005 ;
        RECT 303.300 51.670 303.440 534.635 ;
        RECT 303.240 51.350 303.500 51.670 ;
        RECT 1642.300 51.350 1642.560 51.670 ;
        RECT 1642.360 17.410 1642.500 51.350 ;
        RECT 1642.360 17.270 1644.340 17.410 ;
        RECT 1644.200 2.400 1644.340 17.270 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
      LAYER via2 ;
        RECT 303.230 534.680 303.510 534.960 ;
      LAYER met3 ;
        RECT 303.205 534.970 303.535 534.985 ;
        RECT 303.205 534.880 310.500 534.970 ;
        RECT 303.205 534.670 314.000 534.880 ;
        RECT 303.205 534.655 303.535 534.670 ;
        RECT 310.000 534.280 314.000 534.670 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1318.430 1336.100 1318.750 1336.160 ;
        RECT 1439.410 1336.100 1439.730 1336.160 ;
        RECT 1318.430 1335.960 1439.730 1336.100 ;
        RECT 1318.430 1335.900 1318.750 1335.960 ;
        RECT 1439.410 1335.900 1439.730 1335.960 ;
        RECT 1439.410 431.360 1439.730 431.420 ;
        RECT 1656.530 431.360 1656.850 431.420 ;
        RECT 1439.410 431.220 1656.850 431.360 ;
        RECT 1439.410 431.160 1439.730 431.220 ;
        RECT 1656.530 431.160 1656.850 431.220 ;
      LAYER via ;
        RECT 1318.460 1335.900 1318.720 1336.160 ;
        RECT 1439.440 1335.900 1439.700 1336.160 ;
        RECT 1439.440 431.160 1439.700 431.420 ;
        RECT 1656.560 431.160 1656.820 431.420 ;
      LAYER met2 ;
        RECT 1318.460 1335.870 1318.720 1336.190 ;
        RECT 1439.440 1335.870 1439.700 1336.190 ;
        RECT 1318.520 1325.025 1318.660 1335.870 ;
        RECT 1318.410 1321.025 1318.690 1325.025 ;
        RECT 1439.500 431.450 1439.640 1335.870 ;
        RECT 1439.440 431.130 1439.700 431.450 ;
        RECT 1656.560 431.130 1656.820 431.450 ;
        RECT 1656.620 17.410 1656.760 431.130 ;
        RECT 1656.620 17.270 1662.280 17.410 ;
        RECT 1662.140 2.400 1662.280 17.270 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1027.710 53.620 1028.030 53.680 ;
        RECT 1676.770 53.620 1677.090 53.680 ;
        RECT 1027.710 53.480 1677.090 53.620 ;
        RECT 1027.710 53.420 1028.030 53.480 ;
        RECT 1676.770 53.420 1677.090 53.480 ;
      LAYER via ;
        RECT 1027.740 53.420 1028.000 53.680 ;
        RECT 1676.800 53.420 1677.060 53.680 ;
      LAYER met2 ;
        RECT 1024.930 216.650 1025.210 220.000 ;
        RECT 1024.930 216.510 1027.940 216.650 ;
        RECT 1024.930 216.000 1025.210 216.510 ;
        RECT 1027.800 53.710 1027.940 216.510 ;
        RECT 1027.740 53.390 1028.000 53.710 ;
        RECT 1676.800 53.390 1677.060 53.710 ;
        RECT 1676.860 17.410 1677.000 53.390 ;
        RECT 1676.860 17.270 1679.760 17.410 ;
        RECT 1679.620 2.400 1679.760 17.270 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1404.910 189.960 1405.230 190.020 ;
        RECT 1697.470 189.960 1697.790 190.020 ;
        RECT 1404.910 189.820 1697.790 189.960 ;
        RECT 1404.910 189.760 1405.230 189.820 ;
        RECT 1697.470 189.760 1697.790 189.820 ;
      LAYER via ;
        RECT 1404.940 189.760 1405.200 190.020 ;
        RECT 1697.500 189.760 1697.760 190.020 ;
      LAYER met2 ;
        RECT 1404.890 216.000 1405.170 220.000 ;
        RECT 1405.000 190.050 1405.140 216.000 ;
        RECT 1404.940 189.730 1405.200 190.050 ;
        RECT 1697.500 189.730 1697.760 190.050 ;
        RECT 1697.560 2.400 1697.700 189.730 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.690 1321.650 314.970 1325.025 ;
        RECT 316.110 1321.650 316.390 1321.765 ;
        RECT 314.690 1321.510 316.390 1321.650 ;
        RECT 314.690 1321.025 314.970 1321.510 ;
        RECT 316.110 1321.395 316.390 1321.510 ;
        RECT 731.490 140.915 731.770 141.285 ;
        RECT 731.560 16.730 731.700 140.915 ;
        RECT 731.560 16.590 734.460 16.730 ;
        RECT 734.320 2.400 734.460 16.590 ;
        RECT 734.110 -4.800 734.670 2.400 ;
      LAYER via2 ;
        RECT 316.110 1321.440 316.390 1321.720 ;
        RECT 731.490 140.960 731.770 141.240 ;
      LAYER met3 ;
        RECT 316.085 1321.730 316.415 1321.745 ;
        RECT 322.270 1321.730 322.650 1321.740 ;
        RECT 316.085 1321.430 322.650 1321.730 ;
        RECT 316.085 1321.415 316.415 1321.430 ;
        RECT 322.270 1321.420 322.650 1321.430 ;
        RECT 322.270 141.250 322.650 141.260 ;
        RECT 731.465 141.250 731.795 141.265 ;
        RECT 322.270 140.950 731.795 141.250 ;
        RECT 322.270 140.940 322.650 140.950 ;
        RECT 731.465 140.935 731.795 140.950 ;
      LAYER via3 ;
        RECT 322.300 1321.420 322.620 1321.740 ;
        RECT 322.300 140.940 322.620 141.260 ;
      LAYER met4 ;
        RECT 322.295 1321.415 322.625 1321.745 ;
        RECT 322.310 141.265 322.610 1321.415 ;
        RECT 322.295 140.935 322.625 141.265 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 862.110 53.280 862.430 53.340 ;
        RECT 1711.270 53.280 1711.590 53.340 ;
        RECT 862.110 53.140 1711.590 53.280 ;
        RECT 862.110 53.080 862.430 53.140 ;
        RECT 1711.270 53.080 1711.590 53.140 ;
      LAYER via ;
        RECT 862.140 53.080 862.400 53.340 ;
        RECT 1711.300 53.080 1711.560 53.340 ;
      LAYER met2 ;
        RECT 861.170 216.650 861.450 220.000 ;
        RECT 861.170 216.510 862.340 216.650 ;
        RECT 861.170 216.000 861.450 216.510 ;
        RECT 862.200 53.370 862.340 216.510 ;
        RECT 862.140 53.050 862.400 53.370 ;
        RECT 1711.300 53.050 1711.560 53.370 ;
        RECT 1711.360 17.410 1711.500 53.050 ;
        RECT 1711.360 17.270 1715.640 17.410 ;
        RECT 1715.500 2.400 1715.640 17.270 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 311.490 176.020 311.810 176.080 ;
        RECT 1731.970 176.020 1732.290 176.080 ;
        RECT 311.490 175.880 1732.290 176.020 ;
        RECT 311.490 175.820 311.810 175.880 ;
        RECT 1731.970 175.820 1732.290 175.880 ;
      LAYER via ;
        RECT 311.520 175.820 311.780 176.080 ;
        RECT 1732.000 175.820 1732.260 176.080 ;
      LAYER met2 ;
        RECT 311.510 269.435 311.790 269.805 ;
        RECT 311.580 176.110 311.720 269.435 ;
        RECT 311.520 175.790 311.780 176.110 ;
        RECT 1732.000 175.790 1732.260 176.110 ;
        RECT 1732.060 17.410 1732.200 175.790 ;
        RECT 1732.060 17.270 1733.580 17.410 ;
        RECT 1733.440 2.400 1733.580 17.270 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
      LAYER via2 ;
        RECT 311.510 269.480 311.790 269.760 ;
      LAYER met3 ;
        RECT 310.000 270.440 314.000 271.040 ;
        RECT 311.270 269.785 311.570 270.440 ;
        RECT 311.270 269.470 311.815 269.785 ;
        RECT 311.485 269.455 311.815 269.470 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 778.850 52.260 779.170 52.320 ;
        RECT 1745.770 52.260 1746.090 52.320 ;
        RECT 778.850 52.120 1746.090 52.260 ;
        RECT 778.850 52.060 779.170 52.120 ;
        RECT 1745.770 52.060 1746.090 52.120 ;
      LAYER via ;
        RECT 778.880 52.060 779.140 52.320 ;
        RECT 1745.800 52.060 1746.060 52.320 ;
      LAYER met2 ;
        RECT 777.450 216.650 777.730 220.000 ;
        RECT 777.450 216.510 779.080 216.650 ;
        RECT 777.450 216.000 777.730 216.510 ;
        RECT 778.940 52.350 779.080 216.510 ;
        RECT 778.880 52.030 779.140 52.350 ;
        RECT 1745.800 52.030 1746.060 52.350 ;
        RECT 1745.860 17.410 1746.000 52.030 ;
        RECT 1745.860 17.270 1751.520 17.410 ;
        RECT 1751.380 2.400 1751.520 17.270 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 851.070 200.500 851.390 200.560 ;
        RECT 855.210 200.500 855.530 200.560 ;
        RECT 851.070 200.360 855.530 200.500 ;
        RECT 851.070 200.300 851.390 200.360 ;
        RECT 855.210 200.300 855.530 200.360 ;
        RECT 855.210 52.600 855.530 52.660 ;
        RECT 1766.470 52.600 1766.790 52.660 ;
        RECT 855.210 52.460 1766.790 52.600 ;
        RECT 855.210 52.400 855.530 52.460 ;
        RECT 1766.470 52.400 1766.790 52.460 ;
      LAYER via ;
        RECT 851.100 200.300 851.360 200.560 ;
        RECT 855.240 200.300 855.500 200.560 ;
        RECT 855.240 52.400 855.500 52.660 ;
        RECT 1766.500 52.400 1766.760 52.660 ;
      LAYER met2 ;
        RECT 851.050 216.000 851.330 220.000 ;
        RECT 851.160 200.590 851.300 216.000 ;
        RECT 851.100 200.270 851.360 200.590 ;
        RECT 855.240 200.270 855.500 200.590 ;
        RECT 855.300 52.690 855.440 200.270 ;
        RECT 855.240 52.370 855.500 52.690 ;
        RECT 1766.500 52.370 1766.760 52.690 ;
        RECT 1766.560 17.410 1766.700 52.370 ;
        RECT 1766.560 17.270 1769.000 17.410 ;
        RECT 1768.860 2.400 1769.000 17.270 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.470 200.500 455.790 200.560 ;
        RECT 461.450 200.500 461.770 200.560 ;
        RECT 455.470 200.360 461.770 200.500 ;
        RECT 455.470 200.300 455.790 200.360 ;
        RECT 461.450 200.300 461.770 200.360 ;
        RECT 461.450 51.920 461.770 51.980 ;
        RECT 1780.730 51.920 1781.050 51.980 ;
        RECT 461.450 51.780 1781.050 51.920 ;
        RECT 461.450 51.720 461.770 51.780 ;
        RECT 1780.730 51.720 1781.050 51.780 ;
        RECT 1780.730 19.620 1781.050 19.680 ;
        RECT 1786.710 19.620 1787.030 19.680 ;
        RECT 1780.730 19.480 1787.030 19.620 ;
        RECT 1780.730 19.420 1781.050 19.480 ;
        RECT 1786.710 19.420 1787.030 19.480 ;
      LAYER via ;
        RECT 455.500 200.300 455.760 200.560 ;
        RECT 461.480 200.300 461.740 200.560 ;
        RECT 461.480 51.720 461.740 51.980 ;
        RECT 1780.760 51.720 1781.020 51.980 ;
        RECT 1780.760 19.420 1781.020 19.680 ;
        RECT 1786.740 19.420 1787.000 19.680 ;
      LAYER met2 ;
        RECT 455.450 216.000 455.730 220.000 ;
        RECT 455.560 200.590 455.700 216.000 ;
        RECT 455.500 200.270 455.760 200.590 ;
        RECT 461.480 200.270 461.740 200.590 ;
        RECT 461.540 52.010 461.680 200.270 ;
        RECT 461.480 51.690 461.740 52.010 ;
        RECT 1780.760 51.690 1781.020 52.010 ;
        RECT 1780.820 19.710 1780.960 51.690 ;
        RECT 1780.760 19.390 1781.020 19.710 ;
        RECT 1786.740 19.390 1787.000 19.710 ;
        RECT 1786.800 2.400 1786.940 19.390 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1610.990 45.460 1611.310 45.520 ;
        RECT 1804.650 45.460 1804.970 45.520 ;
        RECT 1610.990 45.320 1804.970 45.460 ;
        RECT 1610.990 45.260 1611.310 45.320 ;
        RECT 1804.650 45.260 1804.970 45.320 ;
      LAYER via ;
        RECT 1611.020 45.260 1611.280 45.520 ;
        RECT 1804.680 45.260 1804.940 45.520 ;
      LAYER met2 ;
        RECT 393.850 1335.675 394.130 1336.045 ;
        RECT 1611.010 1335.675 1611.290 1336.045 ;
        RECT 393.920 1325.025 394.060 1335.675 ;
        RECT 393.810 1321.025 394.090 1325.025 ;
        RECT 1611.080 45.550 1611.220 1335.675 ;
        RECT 1611.020 45.230 1611.280 45.550 ;
        RECT 1804.680 45.230 1804.940 45.550 ;
        RECT 1804.740 2.400 1804.880 45.230 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
      LAYER via2 ;
        RECT 393.850 1335.720 394.130 1336.000 ;
        RECT 1611.010 1335.720 1611.290 1336.000 ;
      LAYER met3 ;
        RECT 393.825 1336.010 394.155 1336.025 ;
        RECT 1610.985 1336.010 1611.315 1336.025 ;
        RECT 393.825 1335.710 1611.315 1336.010 ;
        RECT 393.825 1335.695 394.155 1335.710 ;
        RECT 1610.985 1335.695 1611.315 1335.710 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 965.610 52.940 965.930 53.000 ;
        RECT 1821.670 52.940 1821.990 53.000 ;
        RECT 965.610 52.800 1821.990 52.940 ;
        RECT 965.610 52.740 965.930 52.800 ;
        RECT 1821.670 52.740 1821.990 52.800 ;
      LAYER via ;
        RECT 965.640 52.740 965.900 53.000 ;
        RECT 1821.700 52.740 1821.960 53.000 ;
      LAYER met2 ;
        RECT 965.130 216.650 965.410 220.000 ;
        RECT 965.130 216.510 965.840 216.650 ;
        RECT 965.130 216.000 965.410 216.510 ;
        RECT 965.700 53.030 965.840 216.510 ;
        RECT 965.640 52.710 965.900 53.030 ;
        RECT 1821.700 52.710 1821.960 53.030 ;
        RECT 1821.760 17.410 1821.900 52.710 ;
        RECT 1821.760 17.270 1822.820 17.410 ;
        RECT 1822.680 2.400 1822.820 17.270 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 992.750 1334.060 993.070 1334.120 ;
        RECT 1409.970 1334.060 1410.290 1334.120 ;
        RECT 992.750 1333.920 1410.290 1334.060 ;
        RECT 992.750 1333.860 993.070 1333.920 ;
        RECT 1409.970 1333.860 1410.290 1333.920 ;
        RECT 1409.970 1293.600 1410.290 1293.660 ;
        RECT 1835.470 1293.600 1835.790 1293.660 ;
        RECT 1409.970 1293.460 1835.790 1293.600 ;
        RECT 1409.970 1293.400 1410.290 1293.460 ;
        RECT 1835.470 1293.400 1835.790 1293.460 ;
      LAYER via ;
        RECT 992.780 1333.860 993.040 1334.120 ;
        RECT 1410.000 1333.860 1410.260 1334.120 ;
        RECT 1410.000 1293.400 1410.260 1293.660 ;
        RECT 1835.500 1293.400 1835.760 1293.660 ;
      LAYER met2 ;
        RECT 992.780 1333.830 993.040 1334.150 ;
        RECT 1410.000 1333.830 1410.260 1334.150 ;
        RECT 992.840 1325.025 992.980 1333.830 ;
        RECT 992.730 1321.025 993.010 1325.025 ;
        RECT 1410.060 1293.690 1410.200 1333.830 ;
        RECT 1410.000 1293.370 1410.260 1293.690 ;
        RECT 1835.500 1293.370 1835.760 1293.690 ;
        RECT 1835.560 17.410 1835.700 1293.370 ;
        RECT 1835.560 17.270 1840.300 17.410 ;
        RECT 1840.160 2.400 1840.300 17.270 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 703.410 72.660 703.730 72.720 ;
        RECT 1856.170 72.660 1856.490 72.720 ;
        RECT 703.410 72.520 1856.490 72.660 ;
        RECT 703.410 72.460 703.730 72.520 ;
        RECT 1856.170 72.460 1856.490 72.520 ;
      LAYER via ;
        RECT 703.440 72.460 703.700 72.720 ;
        RECT 1856.200 72.460 1856.460 72.720 ;
      LAYER met2 ;
        RECT 702.930 216.650 703.210 220.000 ;
        RECT 702.930 216.510 703.640 216.650 ;
        RECT 702.930 216.000 703.210 216.510 ;
        RECT 703.500 72.750 703.640 216.510 ;
        RECT 703.440 72.430 703.700 72.750 ;
        RECT 1856.200 72.430 1856.460 72.750 ;
        RECT 1856.260 17.410 1856.400 72.430 ;
        RECT 1856.260 17.270 1858.240 17.410 ;
        RECT 1858.100 2.400 1858.240 17.270 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 576.910 1336.100 577.230 1336.160 ;
        RECT 1289.910 1336.100 1290.230 1336.160 ;
        RECT 576.910 1335.960 1290.230 1336.100 ;
        RECT 576.910 1335.900 577.230 1335.960 ;
        RECT 1289.910 1335.900 1290.230 1335.960 ;
        RECT 1289.910 1328.620 1290.230 1328.680 ;
        RECT 1869.970 1328.620 1870.290 1328.680 ;
        RECT 1289.910 1328.480 1870.290 1328.620 ;
        RECT 1289.910 1328.420 1290.230 1328.480 ;
        RECT 1869.970 1328.420 1870.290 1328.480 ;
        RECT 1869.970 16.900 1870.290 16.960 ;
        RECT 1875.950 16.900 1876.270 16.960 ;
        RECT 1869.970 16.760 1876.270 16.900 ;
        RECT 1869.970 16.700 1870.290 16.760 ;
        RECT 1875.950 16.700 1876.270 16.760 ;
      LAYER via ;
        RECT 576.940 1335.900 577.200 1336.160 ;
        RECT 1289.940 1335.900 1290.200 1336.160 ;
        RECT 1289.940 1328.420 1290.200 1328.680 ;
        RECT 1870.000 1328.420 1870.260 1328.680 ;
        RECT 1870.000 16.700 1870.260 16.960 ;
        RECT 1875.980 16.700 1876.240 16.960 ;
      LAYER met2 ;
        RECT 576.940 1335.870 577.200 1336.190 ;
        RECT 1289.940 1335.870 1290.200 1336.190 ;
        RECT 577.000 1325.025 577.140 1335.870 ;
        RECT 1290.000 1328.710 1290.140 1335.870 ;
        RECT 1289.940 1328.390 1290.200 1328.710 ;
        RECT 1870.000 1328.390 1870.260 1328.710 ;
        RECT 576.890 1321.025 577.170 1325.025 ;
        RECT 1870.060 16.990 1870.200 1328.390 ;
        RECT 1870.000 16.670 1870.260 16.990 ;
        RECT 1875.980 16.670 1876.240 16.990 ;
        RECT 1876.040 2.400 1876.180 16.670 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 311.105 338.045 311.275 386.155 ;
        RECT 448.645 16.745 448.815 17.595 ;
        RECT 507.065 16.065 507.235 17.595 ;
        RECT 531.445 14.365 531.615 16.235 ;
        RECT 568.705 14.365 568.875 15.215 ;
      LAYER mcon ;
        RECT 311.105 385.985 311.275 386.155 ;
        RECT 448.645 17.425 448.815 17.595 ;
        RECT 507.065 17.425 507.235 17.595 ;
        RECT 531.445 16.065 531.615 16.235 ;
        RECT 568.705 15.045 568.875 15.215 ;
      LAYER met1 ;
        RECT 300.450 494.600 300.770 494.660 ;
        RECT 311.490 494.600 311.810 494.660 ;
        RECT 300.450 494.460 311.810 494.600 ;
        RECT 300.450 494.400 300.770 494.460 ;
        RECT 311.490 494.400 311.810 494.460 ;
        RECT 311.030 386.140 311.350 386.200 ;
        RECT 310.835 386.000 311.350 386.140 ;
        RECT 311.030 385.940 311.350 386.000 ;
        RECT 311.045 338.200 311.335 338.245 ;
        RECT 311.490 338.200 311.810 338.260 ;
        RECT 311.045 338.060 311.810 338.200 ;
        RECT 311.045 338.015 311.335 338.060 ;
        RECT 311.490 338.000 311.810 338.060 ;
        RECT 448.585 17.580 448.875 17.625 ;
        RECT 507.005 17.580 507.295 17.625 ;
        RECT 448.585 17.440 507.295 17.580 ;
        RECT 448.585 17.395 448.875 17.440 ;
        RECT 507.005 17.395 507.295 17.440 ;
        RECT 312.410 16.900 312.730 16.960 ;
        RECT 448.585 16.900 448.875 16.945 ;
        RECT 312.410 16.760 448.875 16.900 ;
        RECT 312.410 16.700 312.730 16.760 ;
        RECT 448.585 16.715 448.875 16.760 ;
        RECT 613.710 16.900 614.030 16.960 ;
        RECT 613.710 16.760 650.740 16.900 ;
        RECT 613.710 16.700 614.030 16.760 ;
        RECT 650.600 16.560 650.740 16.760 ;
        RECT 752.170 16.560 752.490 16.620 ;
        RECT 650.600 16.420 752.490 16.560 ;
        RECT 752.170 16.360 752.490 16.420 ;
        RECT 507.005 16.220 507.295 16.265 ;
        RECT 531.385 16.220 531.675 16.265 ;
        RECT 507.005 16.080 531.675 16.220 ;
        RECT 507.005 16.035 507.295 16.080 ;
        RECT 531.385 16.035 531.675 16.080 ;
        RECT 568.645 15.200 568.935 15.245 ;
        RECT 613.710 15.200 614.030 15.260 ;
        RECT 568.645 15.060 614.030 15.200 ;
        RECT 568.645 15.015 568.935 15.060 ;
        RECT 613.710 15.000 614.030 15.060 ;
        RECT 531.385 14.520 531.675 14.565 ;
        RECT 568.645 14.520 568.935 14.565 ;
        RECT 531.385 14.380 568.935 14.520 ;
        RECT 531.385 14.335 531.675 14.380 ;
        RECT 568.645 14.335 568.935 14.380 ;
      LAYER via ;
        RECT 300.480 494.400 300.740 494.660 ;
        RECT 311.520 494.400 311.780 494.660 ;
        RECT 311.060 385.940 311.320 386.200 ;
        RECT 311.520 338.000 311.780 338.260 ;
        RECT 312.440 16.700 312.700 16.960 ;
        RECT 613.740 16.700 614.000 16.960 ;
        RECT 752.200 16.360 752.460 16.620 ;
        RECT 613.740 15.000 614.000 15.260 ;
      LAYER met2 ;
        RECT 300.470 768.555 300.750 768.925 ;
        RECT 300.540 494.690 300.680 768.555 ;
        RECT 311.580 494.690 312.640 494.770 ;
        RECT 300.480 494.370 300.740 494.690 ;
        RECT 311.520 494.630 312.640 494.690 ;
        RECT 311.520 494.370 311.780 494.630 ;
        RECT 312.500 424.730 312.640 494.630 ;
        RECT 311.120 424.590 312.640 424.730 ;
        RECT 311.120 386.230 311.260 424.590 ;
        RECT 311.060 385.910 311.320 386.230 ;
        RECT 311.520 337.970 311.780 338.290 ;
        RECT 311.580 279.210 311.720 337.970 ;
        RECT 310.660 279.070 311.720 279.210 ;
        RECT 310.660 175.170 310.800 279.070 ;
        RECT 310.660 175.030 312.640 175.170 ;
        RECT 312.500 16.990 312.640 175.030 ;
        RECT 312.440 16.670 312.700 16.990 ;
        RECT 613.740 16.670 614.000 16.990 ;
        RECT 613.800 15.290 613.940 16.670 ;
        RECT 752.200 16.330 752.460 16.650 ;
        RECT 613.740 14.970 614.000 15.290 ;
        RECT 752.260 2.400 752.400 16.330 ;
        RECT 752.050 -4.800 752.610 2.400 ;
      LAYER via2 ;
        RECT 300.470 768.600 300.750 768.880 ;
      LAYER met3 ;
        RECT 300.445 768.890 300.775 768.905 ;
        RECT 300.445 768.800 310.500 768.890 ;
        RECT 300.445 768.590 314.000 768.800 ;
        RECT 300.445 768.575 300.775 768.590 ;
        RECT 310.000 768.200 314.000 768.590 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.690 148.395 1890.970 148.765 ;
        RECT 1890.760 17.410 1890.900 148.395 ;
        RECT 1890.760 17.270 1894.120 17.410 ;
        RECT 1893.980 2.400 1894.120 17.270 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
      LAYER via2 ;
        RECT 1890.690 148.440 1890.970 148.720 ;
      LAYER met3 ;
        RECT 303.870 1236.730 304.250 1236.740 ;
        RECT 303.870 1236.640 310.500 1236.730 ;
        RECT 303.870 1236.430 314.000 1236.640 ;
        RECT 303.870 1236.420 304.250 1236.430 ;
        RECT 310.000 1236.040 314.000 1236.430 ;
        RECT 303.870 148.730 304.250 148.740 ;
        RECT 1890.665 148.730 1890.995 148.745 ;
        RECT 303.870 148.430 1890.995 148.730 ;
        RECT 303.870 148.420 304.250 148.430 ;
        RECT 1890.665 148.415 1890.995 148.430 ;
      LAYER via3 ;
        RECT 303.900 1236.420 304.220 1236.740 ;
        RECT 303.900 148.420 304.220 148.740 ;
      LAYER met4 ;
        RECT 303.895 1236.415 304.225 1236.745 ;
        RECT 303.910 148.745 304.210 1236.415 ;
        RECT 303.895 148.415 304.225 148.745 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 938.640 1421.330 938.700 ;
        RECT 1824.890 938.640 1825.210 938.700 ;
        RECT 1421.010 938.500 1825.210 938.640 ;
        RECT 1421.010 938.440 1421.330 938.500 ;
        RECT 1824.890 938.440 1825.210 938.500 ;
        RECT 1824.890 51.920 1825.210 51.980 ;
        RECT 1911.370 51.920 1911.690 51.980 ;
        RECT 1824.890 51.780 1911.690 51.920 ;
        RECT 1824.890 51.720 1825.210 51.780 ;
        RECT 1911.370 51.720 1911.690 51.780 ;
      LAYER via ;
        RECT 1421.040 938.440 1421.300 938.700 ;
        RECT 1824.920 938.440 1825.180 938.700 ;
        RECT 1824.920 51.720 1825.180 51.980 ;
        RECT 1911.400 51.720 1911.660 51.980 ;
      LAYER met2 ;
        RECT 1421.030 943.995 1421.310 944.365 ;
        RECT 1421.100 938.730 1421.240 943.995 ;
        RECT 1421.040 938.410 1421.300 938.730 ;
        RECT 1824.920 938.410 1825.180 938.730 ;
        RECT 1824.980 52.010 1825.120 938.410 ;
        RECT 1824.920 51.690 1825.180 52.010 ;
        RECT 1911.400 51.690 1911.660 52.010 ;
        RECT 1911.460 17.410 1911.600 51.690 ;
        RECT 1911.460 17.270 1912.060 17.410 ;
        RECT 1911.920 2.400 1912.060 17.270 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
      LAYER via2 ;
        RECT 1421.030 944.040 1421.310 944.320 ;
      LAYER met3 ;
        RECT 1421.005 944.330 1421.335 944.345 ;
        RECT 1408.060 944.240 1421.335 944.330 ;
        RECT 1404.305 944.030 1421.335 944.240 ;
        RECT 1404.305 943.640 1408.305 944.030 ;
        RECT 1421.005 944.015 1421.335 944.030 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 814.540 1419.490 814.600 ;
        RECT 1859.390 814.540 1859.710 814.600 ;
        RECT 1419.170 814.400 1859.710 814.540 ;
        RECT 1419.170 814.340 1419.490 814.400 ;
        RECT 1859.390 814.340 1859.710 814.400 ;
        RECT 1859.390 52.260 1859.710 52.320 ;
        RECT 1925.170 52.260 1925.490 52.320 ;
        RECT 1859.390 52.120 1925.490 52.260 ;
        RECT 1859.390 52.060 1859.710 52.120 ;
        RECT 1925.170 52.060 1925.490 52.120 ;
      LAYER via ;
        RECT 1419.200 814.340 1419.460 814.600 ;
        RECT 1859.420 814.340 1859.680 814.600 ;
        RECT 1859.420 52.060 1859.680 52.320 ;
        RECT 1925.200 52.060 1925.460 52.320 ;
      LAYER met2 ;
        RECT 1419.190 818.875 1419.470 819.245 ;
        RECT 1419.260 814.630 1419.400 818.875 ;
        RECT 1419.200 814.310 1419.460 814.630 ;
        RECT 1859.420 814.310 1859.680 814.630 ;
        RECT 1859.480 52.350 1859.620 814.310 ;
        RECT 1859.420 52.030 1859.680 52.350 ;
        RECT 1925.200 52.030 1925.460 52.350 ;
        RECT 1925.260 17.410 1925.400 52.030 ;
        RECT 1925.260 17.270 1929.540 17.410 ;
        RECT 1929.400 2.400 1929.540 17.270 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
      LAYER via2 ;
        RECT 1419.190 818.920 1419.470 819.200 ;
      LAYER met3 ;
        RECT 1419.165 819.210 1419.495 819.225 ;
        RECT 1408.060 819.120 1419.495 819.210 ;
        RECT 1404.305 818.910 1419.495 819.120 ;
        RECT 1404.305 818.520 1408.305 818.910 ;
        RECT 1419.165 818.895 1419.495 818.910 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1083.480 1421.330 1083.540 ;
        RECT 1928.390 1083.480 1928.710 1083.540 ;
        RECT 1421.010 1083.340 1928.710 1083.480 ;
        RECT 1421.010 1083.280 1421.330 1083.340 ;
        RECT 1928.390 1083.280 1928.710 1083.340 ;
        RECT 1928.390 54.980 1928.710 55.040 ;
        RECT 1945.870 54.980 1946.190 55.040 ;
        RECT 1928.390 54.840 1946.190 54.980 ;
        RECT 1928.390 54.780 1928.710 54.840 ;
        RECT 1945.870 54.780 1946.190 54.840 ;
      LAYER via ;
        RECT 1421.040 1083.280 1421.300 1083.540 ;
        RECT 1928.420 1083.280 1928.680 1083.540 ;
        RECT 1928.420 54.780 1928.680 55.040 ;
        RECT 1945.900 54.780 1946.160 55.040 ;
      LAYER met2 ;
        RECT 1421.030 1089.515 1421.310 1089.885 ;
        RECT 1421.100 1083.570 1421.240 1089.515 ;
        RECT 1421.040 1083.250 1421.300 1083.570 ;
        RECT 1928.420 1083.250 1928.680 1083.570 ;
        RECT 1928.480 55.070 1928.620 1083.250 ;
        RECT 1928.420 54.750 1928.680 55.070 ;
        RECT 1945.900 54.750 1946.160 55.070 ;
        RECT 1945.960 17.410 1946.100 54.750 ;
        RECT 1945.960 17.270 1947.480 17.410 ;
        RECT 1947.340 2.400 1947.480 17.270 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1089.560 1421.310 1089.840 ;
      LAYER met3 ;
        RECT 1421.005 1089.850 1421.335 1089.865 ;
        RECT 1408.060 1089.760 1421.335 1089.850 ;
        RECT 1404.305 1089.550 1421.335 1089.760 ;
        RECT 1404.305 1089.160 1408.305 1089.550 ;
        RECT 1421.005 1089.535 1421.335 1089.550 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 629.350 200.500 629.670 200.560 ;
        RECT 633.950 200.500 634.270 200.560 ;
        RECT 629.350 200.360 634.270 200.500 ;
        RECT 629.350 200.300 629.670 200.360 ;
        RECT 633.950 200.300 634.270 200.360 ;
        RECT 633.950 127.740 634.270 127.800 ;
        RECT 1959.670 127.740 1959.990 127.800 ;
        RECT 633.950 127.600 1959.990 127.740 ;
        RECT 633.950 127.540 634.270 127.600 ;
        RECT 1959.670 127.540 1959.990 127.600 ;
      LAYER via ;
        RECT 629.380 200.300 629.640 200.560 ;
        RECT 633.980 200.300 634.240 200.560 ;
        RECT 633.980 127.540 634.240 127.800 ;
        RECT 1959.700 127.540 1959.960 127.800 ;
      LAYER met2 ;
        RECT 629.330 216.000 629.610 220.000 ;
        RECT 629.440 200.590 629.580 216.000 ;
        RECT 629.380 200.270 629.640 200.590 ;
        RECT 633.980 200.270 634.240 200.590 ;
        RECT 634.040 127.830 634.180 200.270 ;
        RECT 633.980 127.510 634.240 127.830 ;
        RECT 1959.700 127.510 1959.960 127.830 ;
        RECT 1959.760 17.410 1959.900 127.510 ;
        RECT 1959.760 17.270 1965.420 17.410 ;
        RECT 1965.280 2.400 1965.420 17.270 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 972.510 1333.720 972.830 1333.780 ;
        RECT 1412.270 1333.720 1412.590 1333.780 ;
        RECT 972.510 1333.580 1412.590 1333.720 ;
        RECT 972.510 1333.520 972.830 1333.580 ;
        RECT 1412.270 1333.520 1412.590 1333.580 ;
        RECT 1410.890 1317.400 1411.210 1317.460 ;
        RECT 1412.270 1317.400 1412.590 1317.460 ;
        RECT 1410.890 1317.260 1412.590 1317.400 ;
        RECT 1410.890 1317.200 1411.210 1317.260 ;
        RECT 1412.270 1317.200 1412.590 1317.260 ;
        RECT 1410.890 1190.240 1411.210 1190.300 ;
        RECT 1980.370 1190.240 1980.690 1190.300 ;
        RECT 1410.890 1190.100 1980.690 1190.240 ;
        RECT 1410.890 1190.040 1411.210 1190.100 ;
        RECT 1980.370 1190.040 1980.690 1190.100 ;
        RECT 1980.370 2.960 1980.690 3.020 ;
        RECT 1983.130 2.960 1983.450 3.020 ;
        RECT 1980.370 2.820 1983.450 2.960 ;
        RECT 1980.370 2.760 1980.690 2.820 ;
        RECT 1983.130 2.760 1983.450 2.820 ;
      LAYER via ;
        RECT 972.540 1333.520 972.800 1333.780 ;
        RECT 1412.300 1333.520 1412.560 1333.780 ;
        RECT 1410.920 1317.200 1411.180 1317.460 ;
        RECT 1412.300 1317.200 1412.560 1317.460 ;
        RECT 1410.920 1190.040 1411.180 1190.300 ;
        RECT 1980.400 1190.040 1980.660 1190.300 ;
        RECT 1980.400 2.760 1980.660 3.020 ;
        RECT 1983.160 2.760 1983.420 3.020 ;
      LAYER met2 ;
        RECT 972.540 1333.490 972.800 1333.810 ;
        RECT 1412.300 1333.490 1412.560 1333.810 ;
        RECT 972.600 1325.025 972.740 1333.490 ;
        RECT 972.490 1321.025 972.770 1325.025 ;
        RECT 1412.360 1317.490 1412.500 1333.490 ;
        RECT 1410.920 1317.170 1411.180 1317.490 ;
        RECT 1412.300 1317.170 1412.560 1317.490 ;
        RECT 1410.980 1190.330 1411.120 1317.170 ;
        RECT 1410.920 1190.010 1411.180 1190.330 ;
        RECT 1980.400 1190.010 1980.660 1190.330 ;
        RECT 1980.460 3.050 1980.600 1190.010 ;
        RECT 1980.400 2.730 1980.660 3.050 ;
        RECT 1983.160 2.730 1983.420 3.050 ;
        RECT 1983.220 2.400 1983.360 2.730 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1439.870 1217.780 1440.190 1217.840 ;
        RECT 2001.070 1217.780 2001.390 1217.840 ;
        RECT 1439.870 1217.640 2001.390 1217.780 ;
        RECT 1439.870 1217.580 1440.190 1217.640 ;
        RECT 2001.070 1217.580 2001.390 1217.640 ;
      LAYER via ;
        RECT 1439.900 1217.580 1440.160 1217.840 ;
        RECT 2001.100 1217.580 2001.360 1217.840 ;
      LAYER met2 ;
        RECT 745.290 1334.315 745.570 1334.685 ;
        RECT 1439.890 1334.315 1440.170 1334.685 ;
        RECT 745.360 1325.025 745.500 1334.315 ;
        RECT 745.250 1321.025 745.530 1325.025 ;
        RECT 1439.960 1217.870 1440.100 1334.315 ;
        RECT 1439.900 1217.550 1440.160 1217.870 ;
        RECT 2001.100 1217.550 2001.360 1217.870 ;
        RECT 2001.160 2.400 2001.300 1217.550 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
      LAYER via2 ;
        RECT 745.290 1334.360 745.570 1334.640 ;
        RECT 1439.890 1334.360 1440.170 1334.640 ;
      LAYER met3 ;
        RECT 745.265 1334.650 745.595 1334.665 ;
        RECT 1439.865 1334.650 1440.195 1334.665 ;
        RECT 745.265 1334.350 1440.195 1334.650 ;
        RECT 745.265 1334.335 745.595 1334.350 ;
        RECT 1439.865 1334.335 1440.195 1334.350 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1353.390 1332.700 1353.710 1332.760 ;
        RECT 1417.790 1332.700 1418.110 1332.760 ;
        RECT 1353.390 1332.560 1418.110 1332.700 ;
        RECT 1353.390 1332.500 1353.710 1332.560 ;
        RECT 1417.790 1332.500 1418.110 1332.560 ;
        RECT 1417.790 1280.000 1418.110 1280.060 ;
        RECT 2014.870 1280.000 2015.190 1280.060 ;
        RECT 1417.790 1279.860 2015.190 1280.000 ;
        RECT 1417.790 1279.800 1418.110 1279.860 ;
        RECT 2014.870 1279.800 2015.190 1279.860 ;
      LAYER via ;
        RECT 1353.420 1332.500 1353.680 1332.760 ;
        RECT 1417.820 1332.500 1418.080 1332.760 ;
        RECT 1417.820 1279.800 1418.080 1280.060 ;
        RECT 2014.900 1279.800 2015.160 1280.060 ;
      LAYER met2 ;
        RECT 1353.420 1332.470 1353.680 1332.790 ;
        RECT 1417.820 1332.470 1418.080 1332.790 ;
        RECT 1353.480 1325.025 1353.620 1332.470 ;
        RECT 1353.370 1321.025 1353.650 1325.025 ;
        RECT 1417.880 1280.090 1418.020 1332.470 ;
        RECT 1417.820 1279.770 1418.080 1280.090 ;
        RECT 2014.900 1279.770 2015.160 1280.090 ;
        RECT 2014.960 16.730 2015.100 1279.770 ;
        RECT 2014.960 16.590 2018.780 16.730 ;
        RECT 2018.640 2.400 2018.780 16.590 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 476.240 1419.490 476.300 ;
        RECT 1949.090 476.240 1949.410 476.300 ;
        RECT 1419.170 476.100 1949.410 476.240 ;
        RECT 1419.170 476.040 1419.490 476.100 ;
        RECT 1949.090 476.040 1949.410 476.100 ;
        RECT 1949.090 51.920 1949.410 51.980 ;
        RECT 2035.570 51.920 2035.890 51.980 ;
        RECT 1949.090 51.780 2035.890 51.920 ;
        RECT 1949.090 51.720 1949.410 51.780 ;
        RECT 2035.570 51.720 2035.890 51.780 ;
      LAYER via ;
        RECT 1419.200 476.040 1419.460 476.300 ;
        RECT 1949.120 476.040 1949.380 476.300 ;
        RECT 1949.120 51.720 1949.380 51.980 ;
        RECT 2035.600 51.720 2035.860 51.980 ;
      LAYER met2 ;
        RECT 1419.190 476.155 1419.470 476.525 ;
        RECT 1419.200 476.010 1419.460 476.155 ;
        RECT 1949.120 476.010 1949.380 476.330 ;
        RECT 1949.180 52.010 1949.320 476.010 ;
        RECT 1949.120 51.690 1949.380 52.010 ;
        RECT 2035.600 51.690 2035.860 52.010 ;
        RECT 2035.660 16.730 2035.800 51.690 ;
        RECT 2035.660 16.590 2036.720 16.730 ;
        RECT 2036.580 2.400 2036.720 16.590 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
      LAYER via2 ;
        RECT 1419.190 476.200 1419.470 476.480 ;
      LAYER met3 ;
        RECT 1419.165 476.490 1419.495 476.505 ;
        RECT 1408.060 476.400 1419.495 476.490 ;
        RECT 1404.305 476.190 1419.495 476.400 ;
        RECT 1404.305 475.800 1408.305 476.190 ;
        RECT 1419.165 476.175 1419.495 476.190 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1419.170 490.180 1419.490 490.240 ;
        RECT 2045.690 490.180 2046.010 490.240 ;
        RECT 1419.170 490.040 2046.010 490.180 ;
        RECT 1419.170 489.980 1419.490 490.040 ;
        RECT 2045.690 489.980 2046.010 490.040 ;
        RECT 2045.690 54.980 2046.010 55.040 ;
        RECT 2049.370 54.980 2049.690 55.040 ;
        RECT 2045.690 54.840 2049.690 54.980 ;
        RECT 2045.690 54.780 2046.010 54.840 ;
        RECT 2049.370 54.780 2049.690 54.840 ;
      LAYER via ;
        RECT 1419.200 489.980 1419.460 490.240 ;
        RECT 2045.720 489.980 2045.980 490.240 ;
        RECT 2045.720 54.780 2045.980 55.040 ;
        RECT 2049.400 54.780 2049.660 55.040 ;
      LAYER met2 ;
        RECT 1419.200 490.125 1419.460 490.270 ;
        RECT 1419.190 489.755 1419.470 490.125 ;
        RECT 2045.720 489.950 2045.980 490.270 ;
        RECT 2045.780 55.070 2045.920 489.950 ;
        RECT 2045.720 54.750 2045.980 55.070 ;
        RECT 2049.400 54.750 2049.660 55.070 ;
        RECT 2049.460 16.730 2049.600 54.750 ;
        RECT 2049.460 16.590 2054.660 16.730 ;
        RECT 2054.520 2.400 2054.660 16.590 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
      LAYER via2 ;
        RECT 1419.190 489.800 1419.470 490.080 ;
      LAYER met3 ;
        RECT 1419.165 490.090 1419.495 490.105 ;
        RECT 1408.060 490.000 1419.495 490.090 ;
        RECT 1404.305 489.790 1419.495 490.000 ;
        RECT 1404.305 489.400 1408.305 489.790 ;
        RECT 1419.165 489.775 1419.495 489.790 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 947.670 1349.360 947.990 1349.420 ;
        RECT 1429.750 1349.360 1430.070 1349.420 ;
        RECT 947.670 1349.220 1430.070 1349.360 ;
        RECT 947.670 1349.160 947.990 1349.220 ;
        RECT 1429.750 1349.160 1430.070 1349.220 ;
        RECT 772.410 211.040 772.730 211.100 ;
        RECT 1429.750 211.040 1430.070 211.100 ;
        RECT 772.410 210.900 1430.070 211.040 ;
        RECT 772.410 210.840 772.730 210.900 ;
        RECT 1429.750 210.840 1430.070 210.900 ;
        RECT 769.650 17.240 769.970 17.300 ;
        RECT 772.410 17.240 772.730 17.300 ;
        RECT 769.650 17.100 772.730 17.240 ;
        RECT 769.650 17.040 769.970 17.100 ;
        RECT 772.410 17.040 772.730 17.100 ;
      LAYER via ;
        RECT 947.700 1349.160 947.960 1349.420 ;
        RECT 1429.780 1349.160 1430.040 1349.420 ;
        RECT 772.440 210.840 772.700 211.100 ;
        RECT 1429.780 210.840 1430.040 211.100 ;
        RECT 769.680 17.040 769.940 17.300 ;
        RECT 772.440 17.040 772.700 17.300 ;
      LAYER met2 ;
        RECT 947.700 1349.130 947.960 1349.450 ;
        RECT 1429.780 1349.130 1430.040 1349.450 ;
        RECT 947.760 1325.025 947.900 1349.130 ;
        RECT 947.650 1321.025 947.930 1325.025 ;
        RECT 1429.840 211.130 1429.980 1349.130 ;
        RECT 772.440 210.810 772.700 211.130 ;
        RECT 1429.780 210.810 1430.040 211.130 ;
        RECT 772.500 17.330 772.640 210.810 ;
        RECT 769.680 17.010 769.940 17.330 ;
        RECT 772.440 17.010 772.700 17.330 ;
        RECT 769.740 2.400 769.880 17.010 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.150 200.500 574.470 200.560 ;
        RECT 579.210 200.500 579.530 200.560 ;
        RECT 574.150 200.360 579.530 200.500 ;
        RECT 574.150 200.300 574.470 200.360 ;
        RECT 579.210 200.300 579.530 200.360 ;
        RECT 579.210 79.800 579.530 79.860 ;
        RECT 2070.070 79.800 2070.390 79.860 ;
        RECT 579.210 79.660 2070.390 79.800 ;
        RECT 579.210 79.600 579.530 79.660 ;
        RECT 2070.070 79.600 2070.390 79.660 ;
      LAYER via ;
        RECT 574.180 200.300 574.440 200.560 ;
        RECT 579.240 200.300 579.500 200.560 ;
        RECT 579.240 79.600 579.500 79.860 ;
        RECT 2070.100 79.600 2070.360 79.860 ;
      LAYER met2 ;
        RECT 574.130 216.000 574.410 220.000 ;
        RECT 574.240 200.590 574.380 216.000 ;
        RECT 574.180 200.270 574.440 200.590 ;
        RECT 579.240 200.270 579.500 200.590 ;
        RECT 579.300 79.890 579.440 200.270 ;
        RECT 579.240 79.570 579.500 79.890 ;
        RECT 2070.100 79.570 2070.360 79.890 ;
        RECT 2070.160 3.130 2070.300 79.570 ;
        RECT 2070.160 2.990 2072.600 3.130 ;
        RECT 2072.460 2.400 2072.600 2.990 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1246.670 200.840 1246.990 200.900 ;
        RECT 1279.790 200.840 1280.110 200.900 ;
        RECT 1246.670 200.700 1280.110 200.840 ;
        RECT 1246.670 200.640 1246.990 200.700 ;
        RECT 1279.790 200.640 1280.110 200.700 ;
        RECT 1279.790 19.280 1280.110 19.340 ;
        RECT 2089.850 19.280 2090.170 19.340 ;
        RECT 1279.790 19.140 2090.170 19.280 ;
        RECT 1279.790 19.080 1280.110 19.140 ;
        RECT 2089.850 19.080 2090.170 19.140 ;
      LAYER via ;
        RECT 1246.700 200.640 1246.960 200.900 ;
        RECT 1279.820 200.640 1280.080 200.900 ;
        RECT 1279.820 19.080 1280.080 19.340 ;
        RECT 2089.880 19.080 2090.140 19.340 ;
      LAYER met2 ;
        RECT 1246.650 216.000 1246.930 220.000 ;
        RECT 1246.760 200.930 1246.900 216.000 ;
        RECT 1246.700 200.610 1246.960 200.930 ;
        RECT 1279.820 200.610 1280.080 200.930 ;
        RECT 1279.880 19.370 1280.020 200.610 ;
        RECT 1279.820 19.050 1280.080 19.370 ;
        RECT 2089.880 19.050 2090.140 19.370 ;
        RECT 2089.940 2.400 2090.080 19.050 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1271.510 200.500 1271.830 200.560 ;
        RECT 1276.110 200.500 1276.430 200.560 ;
        RECT 1271.510 200.360 1276.430 200.500 ;
        RECT 1271.510 200.300 1271.830 200.360 ;
        RECT 1276.110 200.300 1276.430 200.360 ;
        RECT 1276.110 18.940 1276.430 19.000 ;
        RECT 2107.790 18.940 2108.110 19.000 ;
        RECT 1276.110 18.800 2108.110 18.940 ;
        RECT 1276.110 18.740 1276.430 18.800 ;
        RECT 2107.790 18.740 2108.110 18.800 ;
      LAYER via ;
        RECT 1271.540 200.300 1271.800 200.560 ;
        RECT 1276.140 200.300 1276.400 200.560 ;
        RECT 1276.140 18.740 1276.400 19.000 ;
        RECT 2107.820 18.740 2108.080 19.000 ;
      LAYER met2 ;
        RECT 1271.490 216.000 1271.770 220.000 ;
        RECT 1271.600 200.590 1271.740 216.000 ;
        RECT 1271.540 200.270 1271.800 200.590 ;
        RECT 1276.140 200.270 1276.400 200.590 ;
        RECT 1276.200 19.030 1276.340 200.270 ;
        RECT 1276.140 18.710 1276.400 19.030 ;
        RECT 2107.820 18.710 2108.080 19.030 ;
        RECT 2107.880 2.400 2108.020 18.710 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 989.990 205.940 990.310 206.000 ;
        RECT 1024.490 205.940 1024.810 206.000 ;
        RECT 989.990 205.800 1024.810 205.940 ;
        RECT 989.990 205.740 990.310 205.800 ;
        RECT 1024.490 205.740 1024.810 205.800 ;
        RECT 1024.490 18.260 1024.810 18.320 ;
        RECT 2125.270 18.260 2125.590 18.320 ;
        RECT 1024.490 18.120 2125.590 18.260 ;
        RECT 1024.490 18.060 1024.810 18.120 ;
        RECT 2125.270 18.060 2125.590 18.120 ;
      LAYER via ;
        RECT 990.020 205.740 990.280 206.000 ;
        RECT 1024.520 205.740 1024.780 206.000 ;
        RECT 1024.520 18.060 1024.780 18.320 ;
        RECT 2125.300 18.060 2125.560 18.320 ;
      LAYER met2 ;
        RECT 989.970 216.000 990.250 220.000 ;
        RECT 990.080 206.030 990.220 216.000 ;
        RECT 990.020 205.710 990.280 206.030 ;
        RECT 1024.520 205.710 1024.780 206.030 ;
        RECT 1024.580 18.350 1024.720 205.710 ;
        RECT 1024.520 18.030 1024.780 18.350 ;
        RECT 2125.300 18.030 2125.560 18.350 ;
        RECT 2125.360 16.730 2125.500 18.030 ;
        RECT 2125.360 16.590 2125.960 16.730 ;
        RECT 2125.820 2.400 2125.960 16.590 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2125.345 16.745 2125.515 17.595 ;
      LAYER mcon ;
        RECT 2125.345 17.425 2125.515 17.595 ;
      LAYER met1 ;
        RECT 415.910 203.900 416.230 203.960 ;
        RECT 575.990 203.900 576.310 203.960 ;
        RECT 415.910 203.760 576.310 203.900 ;
        RECT 415.910 203.700 416.230 203.760 ;
        RECT 575.990 203.700 576.310 203.760 ;
        RECT 575.990 17.580 576.310 17.640 ;
        RECT 2125.285 17.580 2125.575 17.625 ;
        RECT 575.990 17.440 2125.575 17.580 ;
        RECT 575.990 17.380 576.310 17.440 ;
        RECT 2125.285 17.395 2125.575 17.440 ;
        RECT 2125.285 16.900 2125.575 16.945 ;
        RECT 2143.670 16.900 2143.990 16.960 ;
        RECT 2125.285 16.760 2143.990 16.900 ;
        RECT 2125.285 16.715 2125.575 16.760 ;
        RECT 2143.670 16.700 2143.990 16.760 ;
      LAYER via ;
        RECT 415.940 203.700 416.200 203.960 ;
        RECT 576.020 203.700 576.280 203.960 ;
        RECT 576.020 17.380 576.280 17.640 ;
        RECT 2143.700 16.700 2143.960 16.960 ;
      LAYER met2 ;
        RECT 415.890 216.000 416.170 220.000 ;
        RECT 416.000 203.990 416.140 216.000 ;
        RECT 415.940 203.670 416.200 203.990 ;
        RECT 576.020 203.670 576.280 203.990 ;
        RECT 576.080 17.670 576.220 203.670 ;
        RECT 576.020 17.350 576.280 17.670 ;
        RECT 2143.700 16.670 2143.960 16.990 ;
        RECT 2143.760 2.400 2143.900 16.670 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2048.985 19.465 2049.155 20.315 ;
      LAYER mcon ;
        RECT 2048.985 20.145 2049.155 20.315 ;
      LAYER met1 ;
        RECT 1421.010 393.620 1421.330 393.680 ;
        RECT 2018.090 393.620 2018.410 393.680 ;
        RECT 1421.010 393.480 2018.410 393.620 ;
        RECT 1421.010 393.420 1421.330 393.480 ;
        RECT 2018.090 393.420 2018.410 393.480 ;
        RECT 2018.090 20.300 2018.410 20.360 ;
        RECT 2048.925 20.300 2049.215 20.345 ;
        RECT 2018.090 20.160 2049.215 20.300 ;
        RECT 2018.090 20.100 2018.410 20.160 ;
        RECT 2048.925 20.115 2049.215 20.160 ;
        RECT 2048.925 19.620 2049.215 19.665 ;
        RECT 2161.610 19.620 2161.930 19.680 ;
        RECT 2048.925 19.480 2161.930 19.620 ;
        RECT 2048.925 19.435 2049.215 19.480 ;
        RECT 2161.610 19.420 2161.930 19.480 ;
      LAYER via ;
        RECT 1421.040 393.420 1421.300 393.680 ;
        RECT 2018.120 393.420 2018.380 393.680 ;
        RECT 2018.120 20.100 2018.380 20.360 ;
        RECT 2161.640 19.420 2161.900 19.680 ;
      LAYER met2 ;
        RECT 1421.030 394.555 1421.310 394.925 ;
        RECT 1421.100 393.710 1421.240 394.555 ;
        RECT 1421.040 393.390 1421.300 393.710 ;
        RECT 2018.120 393.390 2018.380 393.710 ;
        RECT 2018.180 20.390 2018.320 393.390 ;
        RECT 2018.120 20.070 2018.380 20.390 ;
        RECT 2161.640 19.390 2161.900 19.710 ;
        RECT 2161.700 2.400 2161.840 19.390 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
      LAYER via2 ;
        RECT 1421.030 394.600 1421.310 394.880 ;
      LAYER met3 ;
        RECT 1421.005 394.890 1421.335 394.905 ;
        RECT 1408.060 394.800 1421.335 394.890 ;
        RECT 1404.305 394.590 1421.335 394.800 ;
        RECT 1404.305 394.200 1408.305 394.590 ;
        RECT 1421.005 394.575 1421.335 394.590 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 821.630 203.900 821.950 203.960 ;
        RECT 2038.790 203.900 2039.110 203.960 ;
        RECT 821.630 203.760 2039.110 203.900 ;
        RECT 821.630 203.700 821.950 203.760 ;
        RECT 2038.790 203.700 2039.110 203.760 ;
        RECT 2038.790 19.960 2039.110 20.020 ;
        RECT 2179.090 19.960 2179.410 20.020 ;
        RECT 2038.790 19.820 2179.410 19.960 ;
        RECT 2038.790 19.760 2039.110 19.820 ;
        RECT 2179.090 19.760 2179.410 19.820 ;
      LAYER via ;
        RECT 821.660 203.700 821.920 203.960 ;
        RECT 2038.820 203.700 2039.080 203.960 ;
        RECT 2038.820 19.760 2039.080 20.020 ;
        RECT 2179.120 19.760 2179.380 20.020 ;
      LAYER met2 ;
        RECT 821.610 216.000 821.890 220.000 ;
        RECT 821.720 203.990 821.860 216.000 ;
        RECT 821.660 203.670 821.920 203.990 ;
        RECT 2038.820 203.670 2039.080 203.990 ;
        RECT 2038.880 20.050 2039.020 203.670 ;
        RECT 2038.820 19.730 2039.080 20.050 ;
        RECT 2179.120 19.730 2179.380 20.050 ;
        RECT 2179.180 2.400 2179.320 19.730 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 295.390 155.280 295.710 155.340 ;
        RECT 2194.270 155.280 2194.590 155.340 ;
        RECT 295.390 155.140 2194.590 155.280 ;
        RECT 295.390 155.080 295.710 155.140 ;
        RECT 2194.270 155.080 2194.590 155.140 ;
      LAYER via ;
        RECT 295.420 155.080 295.680 155.340 ;
        RECT 2194.300 155.080 2194.560 155.340 ;
      LAYER met2 ;
        RECT 295.410 1147.995 295.690 1148.365 ;
        RECT 295.480 155.370 295.620 1147.995 ;
        RECT 295.420 155.050 295.680 155.370 ;
        RECT 2194.300 155.050 2194.560 155.370 ;
        RECT 2194.360 17.410 2194.500 155.050 ;
        RECT 2194.360 17.270 2197.260 17.410 ;
        RECT 2197.120 2.400 2197.260 17.270 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
      LAYER via2 ;
        RECT 295.410 1148.040 295.690 1148.320 ;
      LAYER met3 ;
        RECT 295.385 1148.330 295.715 1148.345 ;
        RECT 295.385 1148.240 310.500 1148.330 ;
        RECT 295.385 1148.030 314.000 1148.240 ;
        RECT 295.385 1148.015 295.715 1148.030 ;
        RECT 310.000 1147.640 314.000 1148.030 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 287.570 876.420 287.890 876.480 ;
        RECT 297.690 876.420 298.010 876.480 ;
        RECT 287.570 876.280 298.010 876.420 ;
        RECT 287.570 876.220 287.890 876.280 ;
        RECT 297.690 876.220 298.010 876.280 ;
        RECT 287.570 86.940 287.890 87.000 ;
        RECT 2215.430 86.940 2215.750 87.000 ;
        RECT 287.570 86.800 2215.750 86.940 ;
        RECT 287.570 86.740 287.890 86.800 ;
        RECT 2215.430 86.740 2215.750 86.800 ;
      LAYER via ;
        RECT 287.600 876.220 287.860 876.480 ;
        RECT 297.720 876.220 297.980 876.480 ;
        RECT 287.600 86.740 287.860 87.000 ;
        RECT 2215.460 86.740 2215.720 87.000 ;
      LAYER met2 ;
        RECT 297.710 877.355 297.990 877.725 ;
        RECT 297.780 876.510 297.920 877.355 ;
        RECT 287.600 876.190 287.860 876.510 ;
        RECT 297.720 876.190 297.980 876.510 ;
        RECT 287.660 87.030 287.800 876.190 ;
        RECT 287.600 86.710 287.860 87.030 ;
        RECT 2215.460 86.710 2215.720 87.030 ;
        RECT 2215.520 7.210 2215.660 86.710 ;
        RECT 2215.060 7.070 2215.660 7.210 ;
        RECT 2215.060 2.400 2215.200 7.070 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
      LAYER via2 ;
        RECT 297.710 877.400 297.990 877.680 ;
      LAYER met3 ;
        RECT 297.685 877.690 298.015 877.705 ;
        RECT 297.685 877.600 310.500 877.690 ;
        RECT 297.685 877.390 314.000 877.600 ;
        RECT 297.685 877.375 298.015 877.390 ;
        RECT 310.000 877.000 314.000 877.390 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1318.045 1314.185 1318.215 1331.695 ;
      LAYER mcon ;
        RECT 1318.045 1331.525 1318.215 1331.695 ;
      LAYER met1 ;
        RECT 1317.970 1331.680 1318.290 1331.740 ;
        RECT 1317.970 1331.540 1318.485 1331.680 ;
        RECT 1317.970 1331.480 1318.290 1331.540 ;
        RECT 1317.985 1314.340 1318.275 1314.385 ;
        RECT 2228.770 1314.340 2229.090 1314.400 ;
        RECT 1317.985 1314.200 2229.090 1314.340 ;
        RECT 1317.985 1314.155 1318.275 1314.200 ;
        RECT 2228.770 1314.140 2229.090 1314.200 ;
      LAYER via ;
        RECT 1318.000 1331.480 1318.260 1331.740 ;
        RECT 2228.800 1314.140 2229.060 1314.400 ;
      LAYER met2 ;
        RECT 710.330 1332.955 710.610 1333.325 ;
        RECT 1317.990 1332.955 1318.270 1333.325 ;
        RECT 710.400 1325.025 710.540 1332.955 ;
        RECT 1318.060 1331.770 1318.200 1332.955 ;
        RECT 1318.000 1331.450 1318.260 1331.770 ;
        RECT 710.290 1321.025 710.570 1325.025 ;
        RECT 2228.800 1314.110 2229.060 1314.430 ;
        RECT 2228.860 17.410 2229.000 1314.110 ;
        RECT 2228.860 17.270 2233.140 17.410 ;
        RECT 2233.000 2.400 2233.140 17.270 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
      LAYER via2 ;
        RECT 710.330 1333.000 710.610 1333.280 ;
        RECT 1317.990 1333.000 1318.270 1333.280 ;
      LAYER met3 ;
        RECT 710.305 1333.290 710.635 1333.305 ;
        RECT 1317.965 1333.290 1318.295 1333.305 ;
        RECT 710.305 1332.990 1318.295 1333.290 ;
        RECT 710.305 1332.975 710.635 1332.990 ;
        RECT 1317.965 1332.975 1318.295 1332.990 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1054.390 206.280 1054.710 206.340 ;
        RECT 1025.040 206.140 1054.710 206.280 ;
        RECT 793.110 205.600 793.430 205.660 ;
        RECT 1025.040 205.600 1025.180 206.140 ;
        RECT 1054.390 206.080 1054.710 206.140 ;
        RECT 793.110 205.460 1025.180 205.600 ;
        RECT 793.110 205.400 793.430 205.460 ;
        RECT 787.590 16.900 787.910 16.960 ;
        RECT 793.110 16.900 793.430 16.960 ;
        RECT 787.590 16.760 793.430 16.900 ;
        RECT 787.590 16.700 787.910 16.760 ;
        RECT 793.110 16.700 793.430 16.760 ;
      LAYER via ;
        RECT 793.140 205.400 793.400 205.660 ;
        RECT 1054.420 206.080 1054.680 206.340 ;
        RECT 787.620 16.700 787.880 16.960 ;
        RECT 793.140 16.700 793.400 16.960 ;
      LAYER met2 ;
        RECT 1054.370 216.000 1054.650 220.000 ;
        RECT 1054.480 206.370 1054.620 216.000 ;
        RECT 1054.420 206.050 1054.680 206.370 ;
        RECT 793.140 205.370 793.400 205.690 ;
        RECT 793.200 16.990 793.340 205.370 ;
        RECT 787.620 16.670 787.880 16.990 ;
        RECT 793.140 16.670 793.400 16.990 ;
        RECT 787.680 2.400 787.820 16.670 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 1325.050 1359.210 1325.165 ;
        RECT 1358.150 1325.025 1359.210 1325.050 ;
        RECT 1357.970 1324.910 1359.210 1325.025 ;
        RECT 1357.970 1321.025 1358.250 1324.910 ;
        RECT 1358.930 1324.795 1359.210 1324.910 ;
        RECT 2250.870 18.515 2251.150 18.885 ;
        RECT 2250.940 2.400 2251.080 18.515 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
      LAYER via2 ;
        RECT 1358.930 1324.840 1359.210 1325.120 ;
        RECT 2250.870 18.560 2251.150 18.840 ;
      LAYER met3 ;
        RECT 1358.905 1325.130 1359.235 1325.145 ;
        RECT 1404.190 1325.130 1404.570 1325.140 ;
        RECT 1358.905 1324.830 1404.570 1325.130 ;
        RECT 1358.905 1324.815 1359.235 1324.830 ;
        RECT 1404.190 1324.820 1404.570 1324.830 ;
        RECT 1404.190 18.850 1404.570 18.860 ;
        RECT 2250.845 18.850 2251.175 18.865 ;
        RECT 1404.190 18.550 2251.175 18.850 ;
        RECT 1404.190 18.540 1404.570 18.550 ;
        RECT 2250.845 18.535 2251.175 18.550 ;
      LAYER via3 ;
        RECT 1404.220 1324.820 1404.540 1325.140 ;
        RECT 1404.220 18.540 1404.540 18.860 ;
      LAYER met4 ;
        RECT 1404.215 1324.815 1404.545 1325.145 ;
        RECT 1404.230 18.865 1404.530 1324.815 ;
        RECT 1404.215 18.535 1404.545 18.865 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 544.710 24.380 545.030 24.440 ;
        RECT 2268.330 24.380 2268.650 24.440 ;
        RECT 544.710 24.240 2268.650 24.380 ;
        RECT 544.710 24.180 545.030 24.240 ;
        RECT 2268.330 24.180 2268.650 24.240 ;
      LAYER via ;
        RECT 544.740 24.180 545.000 24.440 ;
        RECT 2268.360 24.180 2268.620 24.440 ;
      LAYER met2 ;
        RECT 544.690 216.000 544.970 220.000 ;
        RECT 544.800 24.470 544.940 216.000 ;
        RECT 544.740 24.150 545.000 24.470 ;
        RECT 2268.360 24.150 2268.620 24.470 ;
        RECT 2268.420 2.400 2268.560 24.150 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.290 1328.195 1205.570 1328.565 ;
        RECT 1205.360 1325.025 1205.500 1328.195 ;
        RECT 1205.250 1321.025 1205.530 1325.025 ;
        RECT 2286.290 17.835 2286.570 18.205 ;
        RECT 2286.360 2.400 2286.500 17.835 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
      LAYER via2 ;
        RECT 1205.290 1328.240 1205.570 1328.520 ;
        RECT 2286.290 17.880 2286.570 18.160 ;
      LAYER met3 ;
        RECT 1205.265 1328.530 1205.595 1328.545 ;
        RECT 1403.270 1328.530 1403.650 1328.540 ;
        RECT 1205.265 1328.230 1403.650 1328.530 ;
        RECT 1205.265 1328.215 1205.595 1328.230 ;
        RECT 1403.270 1328.220 1403.650 1328.230 ;
        RECT 1403.270 18.170 1403.650 18.180 ;
        RECT 2286.265 18.170 2286.595 18.185 ;
        RECT 1403.270 17.870 2286.595 18.170 ;
        RECT 1403.270 17.860 1403.650 17.870 ;
        RECT 2286.265 17.855 2286.595 17.870 ;
      LAYER via3 ;
        RECT 1403.300 1328.220 1403.620 1328.540 ;
        RECT 1403.300 17.860 1403.620 18.180 ;
      LAYER met4 ;
        RECT 1403.295 1328.215 1403.625 1328.545 ;
        RECT 1403.310 18.185 1403.610 1328.215 ;
        RECT 1403.295 17.855 1403.625 18.185 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1421.010 1021.940 1421.330 1022.000 ;
        RECT 1528.190 1021.940 1528.510 1022.000 ;
        RECT 1421.010 1021.800 1528.510 1021.940 ;
        RECT 1421.010 1021.740 1421.330 1021.800 ;
        RECT 1528.190 1021.740 1528.510 1021.800 ;
        RECT 1528.190 251.840 1528.510 251.900 ;
        RECT 2298.230 251.840 2298.550 251.900 ;
        RECT 1528.190 251.700 2298.550 251.840 ;
        RECT 1528.190 251.640 1528.510 251.700 ;
        RECT 2298.230 251.640 2298.550 251.700 ;
        RECT 2298.230 18.260 2298.550 18.320 ;
        RECT 2304.210 18.260 2304.530 18.320 ;
        RECT 2298.230 18.120 2304.530 18.260 ;
        RECT 2298.230 18.060 2298.550 18.120 ;
        RECT 2304.210 18.060 2304.530 18.120 ;
      LAYER via ;
        RECT 1421.040 1021.740 1421.300 1022.000 ;
        RECT 1528.220 1021.740 1528.480 1022.000 ;
        RECT 1528.220 251.640 1528.480 251.900 ;
        RECT 2298.260 251.640 2298.520 251.900 ;
        RECT 2298.260 18.060 2298.520 18.320 ;
        RECT 2304.240 18.060 2304.500 18.320 ;
      LAYER met2 ;
        RECT 1421.030 1024.235 1421.310 1024.605 ;
        RECT 1421.100 1022.030 1421.240 1024.235 ;
        RECT 1421.040 1021.710 1421.300 1022.030 ;
        RECT 1528.220 1021.710 1528.480 1022.030 ;
        RECT 1528.280 251.930 1528.420 1021.710 ;
        RECT 1528.220 251.610 1528.480 251.930 ;
        RECT 2298.260 251.610 2298.520 251.930 ;
        RECT 2298.320 18.350 2298.460 251.610 ;
        RECT 2298.260 18.030 2298.520 18.350 ;
        RECT 2304.240 18.030 2304.500 18.350 ;
        RECT 2304.300 2.400 2304.440 18.030 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
      LAYER via2 ;
        RECT 1421.030 1024.280 1421.310 1024.560 ;
      LAYER met3 ;
        RECT 1421.005 1024.570 1421.335 1024.585 ;
        RECT 1408.060 1024.480 1421.335 1024.570 ;
        RECT 1404.305 1024.270 1421.335 1024.480 ;
        RECT 1404.305 1023.880 1408.305 1024.270 ;
        RECT 1421.005 1024.255 1421.335 1024.270 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1783.490 51.580 1783.810 51.640 ;
        RECT 2318.470 51.580 2318.790 51.640 ;
        RECT 1783.490 51.440 2318.790 51.580 ;
        RECT 1783.490 51.380 1783.810 51.440 ;
        RECT 2318.470 51.380 2318.790 51.440 ;
      LAYER via ;
        RECT 1783.520 51.380 1783.780 51.640 ;
        RECT 2318.500 51.380 2318.760 51.640 ;
      LAYER met2 ;
        RECT 645.930 1332.275 646.210 1332.645 ;
        RECT 1783.510 1332.275 1783.790 1332.645 ;
        RECT 646.000 1325.025 646.140 1332.275 ;
        RECT 645.890 1321.025 646.170 1325.025 ;
        RECT 1783.580 51.670 1783.720 1332.275 ;
        RECT 1783.520 51.350 1783.780 51.670 ;
        RECT 2318.500 51.350 2318.760 51.670 ;
        RECT 2318.560 17.410 2318.700 51.350 ;
        RECT 2318.560 17.270 2322.380 17.410 ;
        RECT 2322.240 2.400 2322.380 17.270 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
      LAYER via2 ;
        RECT 645.930 1332.320 646.210 1332.600 ;
        RECT 1783.510 1332.320 1783.790 1332.600 ;
      LAYER met3 ;
        RECT 645.905 1332.610 646.235 1332.625 ;
        RECT 1783.485 1332.610 1783.815 1332.625 ;
        RECT 645.905 1332.310 1783.815 1332.610 ;
        RECT 645.905 1332.295 646.235 1332.310 ;
        RECT 1783.485 1332.295 1783.815 1332.310 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1249.430 1335.760 1249.750 1335.820 ;
        RECT 1411.350 1335.760 1411.670 1335.820 ;
        RECT 1249.430 1335.620 1411.670 1335.760 ;
        RECT 1249.430 1335.560 1249.750 1335.620 ;
        RECT 1411.350 1335.560 1411.670 1335.620 ;
        RECT 1411.350 1286.800 1411.670 1286.860 ;
        RECT 2339.170 1286.800 2339.490 1286.860 ;
        RECT 1411.350 1286.660 2339.490 1286.800 ;
        RECT 1411.350 1286.600 1411.670 1286.660 ;
        RECT 2339.170 1286.600 2339.490 1286.660 ;
      LAYER via ;
        RECT 1249.460 1335.560 1249.720 1335.820 ;
        RECT 1411.380 1335.560 1411.640 1335.820 ;
        RECT 1411.380 1286.600 1411.640 1286.860 ;
        RECT 2339.200 1286.600 2339.460 1286.860 ;
      LAYER met2 ;
        RECT 1249.460 1335.530 1249.720 1335.850 ;
        RECT 1411.380 1335.530 1411.640 1335.850 ;
        RECT 1249.520 1325.025 1249.660 1335.530 ;
        RECT 1249.410 1321.025 1249.690 1325.025 ;
        RECT 1411.440 1286.890 1411.580 1335.530 ;
        RECT 1411.380 1286.570 1411.640 1286.890 ;
        RECT 2339.200 1286.570 2339.460 1286.890 ;
        RECT 2339.260 7.890 2339.400 1286.570 ;
        RECT 2339.260 7.750 2339.860 7.890 ;
        RECT 2339.720 2.400 2339.860 7.750 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1079.230 200.500 1079.550 200.560 ;
        RECT 1082.910 200.500 1083.230 200.560 ;
        RECT 1079.230 200.360 1083.230 200.500 ;
        RECT 1079.230 200.300 1079.550 200.360 ;
        RECT 1082.910 200.300 1083.230 200.360 ;
        RECT 1082.910 17.920 1083.230 17.980 ;
        RECT 2357.570 17.920 2357.890 17.980 ;
        RECT 1082.910 17.780 2357.890 17.920 ;
        RECT 1082.910 17.720 1083.230 17.780 ;
        RECT 2357.570 17.720 2357.890 17.780 ;
      LAYER via ;
        RECT 1079.260 200.300 1079.520 200.560 ;
        RECT 1082.940 200.300 1083.200 200.560 ;
        RECT 1082.940 17.720 1083.200 17.980 ;
        RECT 2357.600 17.720 2357.860 17.980 ;
      LAYER met2 ;
        RECT 1079.210 216.000 1079.490 220.000 ;
        RECT 1079.320 200.590 1079.460 216.000 ;
        RECT 1079.260 200.270 1079.520 200.590 ;
        RECT 1082.940 200.270 1083.200 200.590 ;
        RECT 1083.000 18.010 1083.140 200.270 ;
        RECT 1082.940 17.690 1083.200 18.010 ;
        RECT 2357.600 17.690 2357.860 18.010 ;
        RECT 2357.660 2.400 2357.800 17.690 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1426.070 18.600 1426.390 18.660 ;
        RECT 2375.510 18.600 2375.830 18.660 ;
        RECT 1426.070 18.460 2375.830 18.600 ;
        RECT 1426.070 18.400 1426.390 18.460 ;
        RECT 2375.510 18.400 2375.830 18.460 ;
      LAYER via ;
        RECT 1426.100 18.400 1426.360 18.660 ;
        RECT 2375.540 18.400 2375.800 18.660 ;
      LAYER met2 ;
        RECT 566.770 1321.650 567.050 1325.025 ;
        RECT 567.730 1321.650 568.010 1321.765 ;
        RECT 566.770 1321.510 568.010 1321.650 ;
        RECT 566.770 1321.025 567.050 1321.510 ;
        RECT 567.730 1321.395 568.010 1321.510 ;
        RECT 1426.090 1319.355 1426.370 1319.725 ;
        RECT 1426.160 18.690 1426.300 1319.355 ;
        RECT 1426.100 18.370 1426.360 18.690 ;
        RECT 2375.540 18.370 2375.800 18.690 ;
        RECT 2375.600 2.400 2375.740 18.370 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
      LAYER via2 ;
        RECT 567.730 1321.440 568.010 1321.720 ;
        RECT 1426.090 1319.400 1426.370 1319.680 ;
      LAYER met3 ;
        RECT 567.705 1321.730 568.035 1321.745 ;
        RECT 567.705 1321.415 568.250 1321.730 ;
        RECT 567.950 1319.690 568.250 1321.415 ;
        RECT 1426.065 1319.690 1426.395 1319.705 ;
        RECT 567.950 1319.390 1426.395 1319.690 ;
        RECT 1426.065 1319.375 1426.395 1319.390 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1148.230 206.280 1148.550 206.340 ;
        RECT 1196.990 206.280 1197.310 206.340 ;
        RECT 1148.230 206.140 1197.310 206.280 ;
        RECT 1148.230 206.080 1148.550 206.140 ;
        RECT 1196.990 206.080 1197.310 206.140 ;
        RECT 1196.990 46.140 1197.310 46.200 ;
        RECT 2393.450 46.140 2393.770 46.200 ;
        RECT 1196.990 46.000 2393.770 46.140 ;
        RECT 1196.990 45.940 1197.310 46.000 ;
        RECT 2393.450 45.940 2393.770 46.000 ;
      LAYER via ;
        RECT 1148.260 206.080 1148.520 206.340 ;
        RECT 1197.020 206.080 1197.280 206.340 ;
        RECT 1197.020 45.940 1197.280 46.200 ;
        RECT 2393.480 45.940 2393.740 46.200 ;
      LAYER met2 ;
        RECT 1148.210 216.000 1148.490 220.000 ;
        RECT 1148.320 206.370 1148.460 216.000 ;
        RECT 1148.260 206.050 1148.520 206.370 ;
        RECT 1197.020 206.050 1197.280 206.370 ;
        RECT 1197.080 46.230 1197.220 206.050 ;
        RECT 1197.020 45.910 1197.280 46.230 ;
        RECT 2393.480 45.910 2393.740 46.230 ;
        RECT 2393.540 2.400 2393.680 45.910 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 748.030 200.500 748.350 200.560 ;
        RECT 751.710 200.500 752.030 200.560 ;
        RECT 748.030 200.360 752.030 200.500 ;
        RECT 748.030 200.300 748.350 200.360 ;
        RECT 751.710 200.300 752.030 200.360 ;
        RECT 2411.390 17.240 2411.710 17.300 ;
        RECT 779.860 17.100 2411.710 17.240 ;
        RECT 751.710 16.900 752.030 16.960 ;
        RECT 779.860 16.900 780.000 17.100 ;
        RECT 2411.390 17.040 2411.710 17.100 ;
        RECT 751.710 16.760 780.000 16.900 ;
        RECT 751.710 16.700 752.030 16.760 ;
      LAYER via ;
        RECT 748.060 200.300 748.320 200.560 ;
        RECT 751.740 200.300 752.000 200.560 ;
        RECT 751.740 16.700 752.000 16.960 ;
        RECT 2411.420 17.040 2411.680 17.300 ;
      LAYER met2 ;
        RECT 748.010 216.000 748.290 220.000 ;
        RECT 748.120 200.590 748.260 216.000 ;
        RECT 748.060 200.270 748.320 200.590 ;
        RECT 751.740 200.270 752.000 200.590 ;
        RECT 751.800 16.990 751.940 200.270 ;
        RECT 2411.420 17.010 2411.680 17.330 ;
        RECT 751.740 16.670 752.000 16.990 ;
        RECT 2411.480 2.400 2411.620 17.010 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 437.145 1318.265 437.315 1321.495 ;
      LAYER mcon ;
        RECT 437.145 1321.325 437.315 1321.495 ;
      LAYER met1 ;
        RECT 437.070 1321.480 437.390 1321.540 ;
        RECT 436.875 1321.340 437.390 1321.480 ;
        RECT 437.070 1321.280 437.390 1321.340 ;
        RECT 275.150 1318.420 275.470 1318.480 ;
        RECT 437.085 1318.420 437.375 1318.465 ;
        RECT 275.150 1318.280 437.375 1318.420 ;
        RECT 275.150 1318.220 275.470 1318.280 ;
        RECT 437.085 1318.235 437.375 1318.280 ;
        RECT 275.150 20.640 275.470 20.700 ;
        RECT 805.530 20.640 805.850 20.700 ;
        RECT 275.150 20.500 805.850 20.640 ;
        RECT 275.150 20.440 275.470 20.500 ;
        RECT 805.530 20.440 805.850 20.500 ;
      LAYER via ;
        RECT 437.100 1321.280 437.360 1321.540 ;
        RECT 275.180 1318.220 275.440 1318.480 ;
        RECT 275.180 20.440 275.440 20.700 ;
        RECT 805.560 20.440 805.820 20.700 ;
      LAYER met2 ;
        RECT 438.890 1321.650 439.170 1325.025 ;
        RECT 437.160 1321.570 439.170 1321.650 ;
        RECT 437.100 1321.510 439.170 1321.570 ;
        RECT 437.100 1321.250 437.360 1321.510 ;
        RECT 438.890 1321.025 439.170 1321.510 ;
        RECT 275.180 1318.190 275.440 1318.510 ;
        RECT 275.240 20.730 275.380 1318.190 ;
        RECT 275.180 20.410 275.440 20.730 ;
        RECT 805.560 20.410 805.820 20.730 ;
        RECT 805.620 2.400 805.760 20.410 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.985 1307.045 25.155 1322.175 ;
        RECT 48.445 1322.005 48.615 1322.855 ;
        RECT 96.285 1321.665 96.455 1322.855 ;
        RECT 145.045 1322.005 145.215 1322.855 ;
        RECT 110.085 1321.665 110.715 1321.835 ;
        RECT 192.885 1321.665 193.055 1322.855 ;
        RECT 207.145 1321.665 207.775 1321.835 ;
        RECT 241.645 1320.645 241.815 1321.835 ;
        RECT 338.245 1320.985 338.415 1321.835 ;
        RECT 362.165 1320.985 362.335 1321.835 ;
        RECT 448.645 1320.645 448.815 1321.495 ;
        RECT 496.485 1321.325 497.115 1321.495 ;
        RECT 531.445 1320.305 531.615 1321.835 ;
        RECT 579.285 1320.305 579.455 1321.155 ;
      LAYER mcon ;
        RECT 48.445 1322.685 48.615 1322.855 ;
        RECT 24.985 1322.005 25.155 1322.175 ;
        RECT 96.285 1322.685 96.455 1322.855 ;
        RECT 145.045 1322.685 145.215 1322.855 ;
        RECT 192.885 1322.685 193.055 1322.855 ;
        RECT 110.545 1321.665 110.715 1321.835 ;
        RECT 207.605 1321.665 207.775 1321.835 ;
        RECT 241.645 1321.665 241.815 1321.835 ;
        RECT 338.245 1321.665 338.415 1321.835 ;
        RECT 362.165 1321.665 362.335 1321.835 ;
        RECT 531.445 1321.665 531.615 1321.835 ;
        RECT 448.645 1321.325 448.815 1321.495 ;
        RECT 496.945 1321.325 497.115 1321.495 ;
        RECT 579.285 1320.985 579.455 1321.155 ;
      LAYER met1 ;
        RECT 664.310 1334.740 664.630 1334.800 ;
        RECT 903.510 1334.740 903.830 1334.800 ;
        RECT 664.310 1334.600 903.830 1334.740 ;
        RECT 664.310 1334.540 664.630 1334.600 ;
        RECT 903.510 1334.540 903.830 1334.600 ;
        RECT 48.385 1322.840 48.675 1322.885 ;
        RECT 96.225 1322.840 96.515 1322.885 ;
        RECT 48.385 1322.700 96.515 1322.840 ;
        RECT 48.385 1322.655 48.675 1322.700 ;
        RECT 96.225 1322.655 96.515 1322.700 ;
        RECT 144.985 1322.840 145.275 1322.885 ;
        RECT 192.825 1322.840 193.115 1322.885 ;
        RECT 144.985 1322.700 193.115 1322.840 ;
        RECT 144.985 1322.655 145.275 1322.700 ;
        RECT 192.825 1322.655 193.115 1322.700 ;
        RECT 24.925 1322.160 25.215 1322.205 ;
        RECT 48.385 1322.160 48.675 1322.205 ;
        RECT 144.985 1322.160 145.275 1322.205 ;
        RECT 664.310 1322.160 664.630 1322.220 ;
        RECT 24.925 1322.020 48.675 1322.160 ;
        RECT 24.925 1321.975 25.215 1322.020 ;
        RECT 48.385 1321.975 48.675 1322.020 ;
        RECT 116.540 1322.020 145.275 1322.160 ;
        RECT 96.225 1321.820 96.515 1321.865 ;
        RECT 110.025 1321.820 110.315 1321.865 ;
        RECT 96.225 1321.680 110.315 1321.820 ;
        RECT 96.225 1321.635 96.515 1321.680 ;
        RECT 110.025 1321.635 110.315 1321.680 ;
        RECT 110.485 1321.820 110.775 1321.865 ;
        RECT 116.540 1321.820 116.680 1322.020 ;
        RECT 144.985 1321.975 145.275 1322.020 ;
        RECT 627.600 1322.020 664.630 1322.160 ;
        RECT 110.485 1321.680 116.680 1321.820 ;
        RECT 192.825 1321.820 193.115 1321.865 ;
        RECT 207.085 1321.820 207.375 1321.865 ;
        RECT 192.825 1321.680 207.375 1321.820 ;
        RECT 110.485 1321.635 110.775 1321.680 ;
        RECT 192.825 1321.635 193.115 1321.680 ;
        RECT 207.085 1321.635 207.375 1321.680 ;
        RECT 207.545 1321.820 207.835 1321.865 ;
        RECT 207.545 1321.680 241.340 1321.820 ;
        RECT 207.545 1321.635 207.835 1321.680 ;
        RECT 241.200 1321.480 241.340 1321.680 ;
        RECT 241.585 1321.635 241.875 1321.865 ;
        RECT 338.185 1321.820 338.475 1321.865 ;
        RECT 362.105 1321.820 362.395 1321.865 ;
        RECT 531.385 1321.820 531.675 1321.865 ;
        RECT 627.600 1321.820 627.740 1322.020 ;
        RECT 664.310 1321.960 664.630 1322.020 ;
        RECT 338.185 1321.680 362.395 1321.820 ;
        RECT 338.185 1321.635 338.475 1321.680 ;
        RECT 362.105 1321.635 362.395 1321.680 ;
        RECT 497.880 1321.680 531.675 1321.820 ;
        RECT 241.660 1321.480 241.800 1321.635 ;
        RECT 241.200 1321.340 241.800 1321.480 ;
        RECT 448.585 1321.480 448.875 1321.525 ;
        RECT 496.425 1321.480 496.715 1321.525 ;
        RECT 448.585 1321.340 496.715 1321.480 ;
        RECT 448.585 1321.295 448.875 1321.340 ;
        RECT 496.425 1321.295 496.715 1321.340 ;
        RECT 496.885 1321.480 497.175 1321.525 ;
        RECT 497.880 1321.480 498.020 1321.680 ;
        RECT 531.385 1321.635 531.675 1321.680 ;
        RECT 592.640 1321.680 627.740 1321.820 ;
        RECT 496.885 1321.340 498.020 1321.480 ;
        RECT 496.885 1321.295 497.175 1321.340 ;
        RECT 338.185 1321.140 338.475 1321.185 ;
        RECT 255.460 1321.000 338.475 1321.140 ;
        RECT 241.585 1320.800 241.875 1320.845 ;
        RECT 255.460 1320.800 255.600 1321.000 ;
        RECT 338.185 1320.955 338.475 1321.000 ;
        RECT 362.105 1321.140 362.395 1321.185 ;
        RECT 579.225 1321.140 579.515 1321.185 ;
        RECT 592.640 1321.140 592.780 1321.680 ;
        RECT 362.105 1321.000 400.500 1321.140 ;
        RECT 362.105 1320.955 362.395 1321.000 ;
        RECT 241.585 1320.660 255.600 1320.800 ;
        RECT 400.360 1320.800 400.500 1321.000 ;
        RECT 579.225 1321.000 592.780 1321.140 ;
        RECT 579.225 1320.955 579.515 1321.000 ;
        RECT 448.585 1320.800 448.875 1320.845 ;
        RECT 400.360 1320.660 448.875 1320.800 ;
        RECT 241.585 1320.615 241.875 1320.660 ;
        RECT 448.585 1320.615 448.875 1320.660 ;
        RECT 531.385 1320.460 531.675 1320.505 ;
        RECT 579.225 1320.460 579.515 1320.505 ;
        RECT 531.385 1320.320 579.515 1320.460 ;
        RECT 531.385 1320.275 531.675 1320.320 ;
        RECT 579.225 1320.275 579.515 1320.320 ;
        RECT 6.510 1307.200 6.830 1307.260 ;
        RECT 24.925 1307.200 25.215 1307.245 ;
        RECT 6.510 1307.060 25.215 1307.200 ;
        RECT 6.510 1307.000 6.830 1307.060 ;
        RECT 24.925 1307.015 25.215 1307.060 ;
        RECT 2.830 17.580 3.150 17.640 ;
        RECT 6.510 17.580 6.830 17.640 ;
        RECT 2.830 17.440 6.830 17.580 ;
        RECT 2.830 17.380 3.150 17.440 ;
        RECT 6.510 17.380 6.830 17.440 ;
      LAYER via ;
        RECT 664.340 1334.540 664.600 1334.800 ;
        RECT 903.540 1334.540 903.800 1334.800 ;
        RECT 664.340 1321.960 664.600 1322.220 ;
        RECT 6.540 1307.000 6.800 1307.260 ;
        RECT 2.860 17.380 3.120 17.640 ;
        RECT 6.540 17.380 6.800 17.640 ;
      LAYER met2 ;
        RECT 664.340 1334.510 664.600 1334.830 ;
        RECT 903.540 1334.510 903.800 1334.830 ;
        RECT 664.400 1322.250 664.540 1334.510 ;
        RECT 903.600 1325.025 903.740 1334.510 ;
        RECT 664.340 1321.930 664.600 1322.250 ;
        RECT 903.490 1321.025 903.770 1325.025 ;
        RECT 6.540 1306.970 6.800 1307.290 ;
        RECT 6.600 17.670 6.740 1306.970 ;
        RECT 2.860 17.350 3.120 17.670 ;
        RECT 6.540 17.350 6.800 17.670 ;
        RECT 2.920 2.400 3.060 17.350 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 13.410 204.580 13.730 204.640 ;
        RECT 1177.670 204.580 1177.990 204.640 ;
        RECT 13.410 204.440 1177.990 204.580 ;
        RECT 13.410 204.380 13.730 204.440 ;
        RECT 1177.670 204.380 1177.990 204.440 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 13.410 17.580 13.730 17.640 ;
        RECT 8.350 17.440 13.730 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 13.410 17.380 13.730 17.440 ;
      LAYER via ;
        RECT 13.440 204.380 13.700 204.640 ;
        RECT 1177.700 204.380 1177.960 204.640 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 13.440 17.380 13.700 17.640 ;
      LAYER met2 ;
        RECT 1177.650 216.000 1177.930 220.000 ;
        RECT 1177.760 204.670 1177.900 216.000 ;
        RECT 13.440 204.350 13.700 204.670 ;
        RECT 1177.700 204.350 1177.960 204.670 ;
        RECT 13.500 17.670 13.640 204.350 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 13.440 17.350 13.700 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 1335.025 367.020 3529.000 ;
        RECT 544.020 1335.025 547.020 3529.000 ;
        RECT 724.020 1335.025 727.020 3529.000 ;
        RECT 904.020 1335.025 907.020 3529.000 ;
        RECT 1084.020 1335.025 1087.020 3529.000 ;
        RECT 1264.020 1335.025 1267.020 3529.000 ;
        RECT 364.020 -9.320 367.020 206.000 ;
        RECT 544.020 -9.320 547.020 206.000 ;
        RECT 724.020 -9.320 727.020 206.000 ;
        RECT 904.020 -9.320 907.020 206.000 ;
        RECT 1084.020 -9.320 1087.020 206.000 ;
        RECT 1264.020 -9.320 1267.020 206.000 ;
        RECT 1444.020 -9.320 1447.020 3529.000 ;
        RECT 1624.020 -9.320 1627.020 3529.000 ;
        RECT 1804.020 -9.320 1807.020 3529.000 ;
        RECT 1984.020 -9.320 1987.020 3529.000 ;
        RECT 2164.020 -9.320 2167.020 3529.000 ;
        RECT 2344.020 -9.320 2347.020 3529.000 ;
        RECT 2524.020 -9.320 2527.020 3529.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 1335.025 457.020 3529.000 ;
        RECT 634.020 1335.025 637.020 3529.000 ;
        RECT 814.020 1335.025 817.020 3529.000 ;
        RECT 994.020 1335.025 997.020 3529.000 ;
        RECT 1174.020 1335.025 1177.020 3529.000 ;
        RECT 1354.020 1335.025 1357.020 3529.000 ;
        RECT 454.020 -9.320 457.020 206.000 ;
        RECT 634.020 -9.320 637.020 206.000 ;
        RECT 814.020 -9.320 817.020 206.000 ;
        RECT 994.020 -9.320 997.020 206.000 ;
        RECT 1174.020 -9.320 1177.020 206.000 ;
        RECT 1354.020 -9.320 1357.020 206.000 ;
        RECT 1534.020 -9.320 1537.020 3529.000 ;
        RECT 1714.020 -9.320 1717.020 3529.000 ;
        RECT 1894.020 -9.320 1897.020 3529.000 ;
        RECT 2074.020 -9.320 2077.020 3529.000 ;
        RECT 2254.020 -9.320 2257.020 3529.000 ;
        RECT 2434.020 -9.320 2437.020 3529.000 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 315.520 226.795 1402.500 1312.245 ;
      LAYER met1 ;
        RECT 312.830 221.820 1403.350 1313.480 ;
      LAYER met2 ;
        RECT 349.650 1321.025 349.930 1325.025 ;
        RECT 354.250 1321.025 354.530 1325.025 ;
        RECT 379.090 1321.025 379.370 1325.025 ;
        RECT 389.210 1321.025 389.490 1325.025 ;
        RECT 403.930 1321.025 404.210 1325.025 ;
        RECT 414.050 1321.025 414.330 1325.025 ;
        RECT 418.650 1321.025 418.930 1325.025 ;
        RECT 453.610 1321.025 453.890 1325.025 ;
        RECT 458.210 1321.025 458.490 1325.025 ;
        RECT 462.810 1321.025 463.090 1325.025 ;
        RECT 468.330 1321.025 468.610 1325.025 ;
        RECT 472.930 1321.025 473.210 1325.025 ;
        RECT 478.450 1321.025 478.730 1325.025 ;
        RECT 502.370 1321.025 502.650 1325.025 ;
        RECT 507.890 1321.025 508.170 1325.025 ;
        RECT 527.210 1321.025 527.490 1325.025 ;
        RECT 547.450 1321.025 547.730 1325.025 ;
        RECT 557.570 1321.025 557.850 1325.025 ;
        RECT 591.610 1321.025 591.890 1325.025 ;
        RECT 597.130 1321.025 597.410 1325.025 ;
        RECT 606.330 1321.025 606.610 1325.025 ;
        RECT 616.450 1321.025 616.730 1325.025 ;
        RECT 626.570 1321.025 626.850 1325.025 ;
        RECT 631.170 1321.025 631.450 1325.025 ;
        RECT 636.690 1321.025 636.970 1325.025 ;
        RECT 651.410 1321.025 651.690 1325.025 ;
        RECT 656.010 1321.025 656.290 1325.025 ;
        RECT 676.250 1321.025 676.530 1325.025 ;
        RECT 690.970 1321.025 691.250 1325.025 ;
        RECT 700.170 1321.025 700.450 1325.025 ;
        RECT 705.690 1321.025 705.970 1325.025 ;
        RECT 730.530 1321.025 730.810 1325.025 ;
        RECT 735.130 1321.025 735.410 1325.025 ;
        RECT 755.370 1321.025 755.650 1325.025 ;
        RECT 759.970 1321.025 760.250 1325.025 ;
        RECT 770.090 1321.025 770.370 1325.025 ;
        RECT 828.970 1321.025 829.250 1325.025 ;
        RECT 834.490 1321.025 834.770 1325.025 ;
        RECT 839.090 1321.025 839.370 1325.025 ;
        RECT 849.210 1321.025 849.490 1325.025 ;
        RECT 878.650 1321.025 878.930 1325.025 ;
        RECT 883.250 1321.025 883.530 1325.025 ;
        RECT 888.770 1321.025 889.050 1325.025 ;
        RECT 913.610 1321.025 913.890 1325.025 ;
        RECT 922.810 1321.025 923.090 1325.025 ;
        RECT 928.330 1321.025 928.610 1325.025 ;
        RECT 932.930 1321.025 933.210 1325.025 ;
        RECT 953.170 1321.025 953.450 1325.025 ;
        RECT 962.370 1321.025 962.650 1325.025 ;
        RECT 967.890 1321.025 968.170 1325.025 ;
        RECT 978.010 1321.025 978.290 1325.025 ;
        RECT 982.610 1321.025 982.890 1325.025 ;
        RECT 1017.570 1321.025 1017.850 1325.025 ;
        RECT 1022.170 1321.025 1022.450 1325.025 ;
        RECT 1026.770 1321.025 1027.050 1325.025 ;
        RECT 1036.890 1321.025 1037.170 1325.025 ;
        RECT 1061.730 1321.025 1062.010 1325.025 ;
        RECT 1086.570 1321.025 1086.850 1325.025 ;
        RECT 1096.690 1321.025 1096.970 1325.025 ;
        RECT 1126.130 1321.025 1126.410 1325.025 ;
        RECT 1136.250 1321.025 1136.530 1325.025 ;
        RECT 1140.850 1321.025 1141.130 1325.025 ;
        RECT 1160.170 1321.025 1160.450 1325.025 ;
        RECT 1170.290 1321.025 1170.570 1325.025 ;
        RECT 1175.810 1321.025 1176.090 1325.025 ;
        RECT 1195.130 1321.025 1195.410 1325.025 ;
        RECT 1199.730 1321.025 1200.010 1325.025 ;
        RECT 1215.370 1321.025 1215.650 1325.025 ;
        RECT 1234.690 1321.025 1234.970 1325.025 ;
        RECT 1239.290 1321.025 1239.570 1325.025 ;
        RECT 1254.930 1321.025 1255.210 1325.025 ;
        RECT 1309.210 1321.025 1309.490 1325.025 ;
        RECT 1334.050 1321.025 1334.330 1325.025 ;
        RECT 1363.490 1321.025 1363.770 1325.025 ;
        RECT 1382.810 1321.025 1383.090 1325.025 ;
      LAYER met2 ;
        RECT 312.860 1320.745 314.410 1321.025 ;
        RECT 315.250 1320.745 319.930 1321.025 ;
        RECT 320.770 1320.745 324.530 1321.025 ;
        RECT 325.370 1320.745 329.130 1321.025 ;
        RECT 329.970 1320.745 334.650 1321.025 ;
        RECT 335.490 1320.745 339.250 1321.025 ;
        RECT 340.090 1320.745 343.850 1321.025 ;
        RECT 344.690 1320.745 349.370 1321.025 ;
        RECT 350.210 1320.745 353.970 1321.025 ;
        RECT 354.810 1320.745 359.490 1321.025 ;
        RECT 360.330 1320.745 364.090 1321.025 ;
        RECT 364.930 1320.745 368.690 1321.025 ;
        RECT 369.530 1320.745 374.210 1321.025 ;
        RECT 375.050 1320.745 378.810 1321.025 ;
        RECT 379.650 1320.745 383.410 1321.025 ;
        RECT 384.250 1320.745 388.930 1321.025 ;
        RECT 389.770 1320.745 393.530 1321.025 ;
        RECT 394.370 1320.745 399.050 1321.025 ;
        RECT 399.890 1320.745 403.650 1321.025 ;
        RECT 404.490 1320.745 408.250 1321.025 ;
        RECT 409.090 1320.745 413.770 1321.025 ;
        RECT 414.610 1320.745 418.370 1321.025 ;
        RECT 419.210 1320.745 422.970 1321.025 ;
        RECT 423.810 1320.745 428.490 1321.025 ;
        RECT 429.330 1320.745 433.090 1321.025 ;
        RECT 433.930 1320.745 438.610 1321.025 ;
        RECT 439.450 1320.745 443.210 1321.025 ;
        RECT 444.050 1320.745 447.810 1321.025 ;
        RECT 448.650 1320.745 453.330 1321.025 ;
        RECT 454.170 1320.745 457.930 1321.025 ;
        RECT 458.770 1320.745 462.530 1321.025 ;
        RECT 463.370 1320.745 468.050 1321.025 ;
        RECT 468.890 1320.745 472.650 1321.025 ;
        RECT 473.490 1320.745 478.170 1321.025 ;
        RECT 479.010 1320.745 482.770 1321.025 ;
        RECT 483.610 1320.745 487.370 1321.025 ;
        RECT 488.210 1320.745 492.890 1321.025 ;
        RECT 493.730 1320.745 497.490 1321.025 ;
        RECT 498.330 1320.745 502.090 1321.025 ;
        RECT 502.930 1320.745 507.610 1321.025 ;
        RECT 508.450 1320.745 512.210 1321.025 ;
        RECT 513.050 1320.745 517.730 1321.025 ;
        RECT 518.570 1320.745 522.330 1321.025 ;
        RECT 523.170 1320.745 526.930 1321.025 ;
        RECT 527.770 1320.745 532.450 1321.025 ;
        RECT 533.290 1320.745 537.050 1321.025 ;
        RECT 537.890 1320.745 541.650 1321.025 ;
        RECT 542.490 1320.745 547.170 1321.025 ;
        RECT 548.010 1320.745 551.770 1321.025 ;
        RECT 552.610 1320.745 557.290 1321.025 ;
        RECT 558.130 1320.745 561.890 1321.025 ;
        RECT 562.730 1320.745 566.490 1321.025 ;
        RECT 567.330 1320.745 572.010 1321.025 ;
        RECT 572.850 1320.745 576.610 1321.025 ;
        RECT 577.450 1320.745 581.210 1321.025 ;
        RECT 582.050 1320.745 586.730 1321.025 ;
        RECT 587.570 1320.745 591.330 1321.025 ;
        RECT 592.170 1320.745 596.850 1321.025 ;
        RECT 597.690 1320.745 601.450 1321.025 ;
        RECT 602.290 1320.745 606.050 1321.025 ;
        RECT 606.890 1320.745 611.570 1321.025 ;
        RECT 612.410 1320.745 616.170 1321.025 ;
        RECT 617.010 1320.745 620.770 1321.025 ;
        RECT 621.610 1320.745 626.290 1321.025 ;
        RECT 627.130 1320.745 630.890 1321.025 ;
        RECT 631.730 1320.745 636.410 1321.025 ;
        RECT 637.250 1320.745 641.010 1321.025 ;
        RECT 641.850 1320.745 645.610 1321.025 ;
        RECT 646.450 1320.745 651.130 1321.025 ;
        RECT 651.970 1320.745 655.730 1321.025 ;
        RECT 656.570 1320.745 660.330 1321.025 ;
        RECT 661.170 1320.745 665.850 1321.025 ;
        RECT 666.690 1320.745 670.450 1321.025 ;
        RECT 671.290 1320.745 675.970 1321.025 ;
        RECT 676.810 1320.745 680.570 1321.025 ;
        RECT 681.410 1320.745 685.170 1321.025 ;
        RECT 686.010 1320.745 690.690 1321.025 ;
        RECT 691.530 1320.745 695.290 1321.025 ;
        RECT 696.130 1320.745 699.890 1321.025 ;
        RECT 700.730 1320.745 705.410 1321.025 ;
        RECT 706.250 1320.745 710.010 1321.025 ;
        RECT 710.850 1320.745 715.530 1321.025 ;
        RECT 716.370 1320.745 720.130 1321.025 ;
        RECT 720.970 1320.745 724.730 1321.025 ;
        RECT 725.570 1320.745 730.250 1321.025 ;
        RECT 731.090 1320.745 734.850 1321.025 ;
        RECT 735.690 1320.745 739.450 1321.025 ;
        RECT 740.290 1320.745 744.970 1321.025 ;
        RECT 745.810 1320.745 749.570 1321.025 ;
        RECT 750.410 1320.745 755.090 1321.025 ;
        RECT 755.930 1320.745 759.690 1321.025 ;
        RECT 760.530 1320.745 764.290 1321.025 ;
        RECT 765.130 1320.745 769.810 1321.025 ;
        RECT 770.650 1320.745 774.410 1321.025 ;
        RECT 775.250 1320.745 779.010 1321.025 ;
        RECT 779.850 1320.745 784.530 1321.025 ;
        RECT 785.370 1320.745 789.130 1321.025 ;
        RECT 789.970 1320.745 794.650 1321.025 ;
        RECT 795.490 1320.745 799.250 1321.025 ;
        RECT 800.090 1320.745 803.850 1321.025 ;
        RECT 804.690 1320.745 809.370 1321.025 ;
        RECT 810.210 1320.745 813.970 1321.025 ;
        RECT 814.810 1320.745 819.490 1321.025 ;
        RECT 820.330 1320.745 824.090 1321.025 ;
        RECT 824.930 1320.745 828.690 1321.025 ;
        RECT 829.530 1320.745 834.210 1321.025 ;
        RECT 835.050 1320.745 838.810 1321.025 ;
        RECT 839.650 1320.745 843.410 1321.025 ;
        RECT 844.250 1320.745 848.930 1321.025 ;
        RECT 849.770 1320.745 853.530 1321.025 ;
        RECT 854.370 1320.745 859.050 1321.025 ;
        RECT 859.890 1320.745 863.650 1321.025 ;
        RECT 864.490 1320.745 868.250 1321.025 ;
        RECT 869.090 1320.745 873.770 1321.025 ;
        RECT 874.610 1320.745 878.370 1321.025 ;
        RECT 879.210 1320.745 882.970 1321.025 ;
        RECT 883.810 1320.745 888.490 1321.025 ;
        RECT 889.330 1320.745 893.090 1321.025 ;
        RECT 893.930 1320.745 898.610 1321.025 ;
        RECT 899.450 1320.745 903.210 1321.025 ;
        RECT 904.050 1320.745 907.810 1321.025 ;
        RECT 908.650 1320.745 913.330 1321.025 ;
        RECT 914.170 1320.745 917.930 1321.025 ;
        RECT 918.770 1320.745 922.530 1321.025 ;
        RECT 923.370 1320.745 928.050 1321.025 ;
        RECT 928.890 1320.745 932.650 1321.025 ;
        RECT 933.490 1320.745 938.170 1321.025 ;
        RECT 939.010 1320.745 942.770 1321.025 ;
        RECT 943.610 1320.745 947.370 1321.025 ;
        RECT 948.210 1320.745 952.890 1321.025 ;
        RECT 953.730 1320.745 957.490 1321.025 ;
        RECT 958.330 1320.745 962.090 1321.025 ;
        RECT 962.930 1320.745 967.610 1321.025 ;
        RECT 968.450 1320.745 972.210 1321.025 ;
        RECT 973.050 1320.745 977.730 1321.025 ;
        RECT 978.570 1320.745 982.330 1321.025 ;
        RECT 983.170 1320.745 986.930 1321.025 ;
        RECT 987.770 1320.745 992.450 1321.025 ;
        RECT 993.290 1320.745 997.050 1321.025 ;
        RECT 997.890 1320.745 1001.650 1321.025 ;
        RECT 1002.490 1320.745 1007.170 1321.025 ;
        RECT 1008.010 1320.745 1011.770 1321.025 ;
        RECT 1012.610 1320.745 1017.290 1321.025 ;
        RECT 1018.130 1320.745 1021.890 1321.025 ;
        RECT 1022.730 1320.745 1026.490 1321.025 ;
        RECT 1027.330 1320.745 1032.010 1321.025 ;
        RECT 1032.850 1320.745 1036.610 1321.025 ;
        RECT 1037.450 1320.745 1041.210 1321.025 ;
        RECT 1042.050 1320.745 1046.730 1321.025 ;
        RECT 1047.570 1320.745 1051.330 1321.025 ;
        RECT 1052.170 1320.745 1056.850 1321.025 ;
        RECT 1057.690 1320.745 1061.450 1321.025 ;
        RECT 1062.290 1320.745 1066.050 1321.025 ;
        RECT 1066.890 1320.745 1071.570 1321.025 ;
        RECT 1072.410 1320.745 1076.170 1321.025 ;
        RECT 1077.010 1320.745 1080.770 1321.025 ;
        RECT 1081.610 1320.745 1086.290 1321.025 ;
        RECT 1087.130 1320.745 1090.890 1321.025 ;
        RECT 1091.730 1320.745 1096.410 1321.025 ;
        RECT 1097.250 1320.745 1101.010 1321.025 ;
        RECT 1101.850 1320.745 1105.610 1321.025 ;
        RECT 1106.450 1320.745 1111.130 1321.025 ;
        RECT 1111.970 1320.745 1115.730 1321.025 ;
        RECT 1116.570 1320.745 1120.330 1321.025 ;
        RECT 1121.170 1320.745 1125.850 1321.025 ;
        RECT 1126.690 1320.745 1130.450 1321.025 ;
        RECT 1131.290 1320.745 1135.970 1321.025 ;
        RECT 1136.810 1320.745 1140.570 1321.025 ;
        RECT 1141.410 1320.745 1145.170 1321.025 ;
        RECT 1146.010 1320.745 1150.690 1321.025 ;
        RECT 1151.530 1320.745 1155.290 1321.025 ;
        RECT 1156.130 1320.745 1159.890 1321.025 ;
        RECT 1160.730 1320.745 1165.410 1321.025 ;
        RECT 1166.250 1320.745 1170.010 1321.025 ;
        RECT 1170.850 1320.745 1175.530 1321.025 ;
        RECT 1176.370 1320.745 1180.130 1321.025 ;
        RECT 1180.970 1320.745 1184.730 1321.025 ;
        RECT 1185.570 1320.745 1190.250 1321.025 ;
        RECT 1191.090 1320.745 1194.850 1321.025 ;
        RECT 1195.690 1320.745 1199.450 1321.025 ;
        RECT 1200.290 1320.745 1204.970 1321.025 ;
        RECT 1205.810 1320.745 1209.570 1321.025 ;
        RECT 1210.410 1320.745 1215.090 1321.025 ;
        RECT 1215.930 1320.745 1219.690 1321.025 ;
        RECT 1220.530 1320.745 1224.290 1321.025 ;
        RECT 1225.130 1320.745 1229.810 1321.025 ;
        RECT 1230.650 1320.745 1234.410 1321.025 ;
        RECT 1235.250 1320.745 1239.010 1321.025 ;
        RECT 1239.850 1320.745 1244.530 1321.025 ;
        RECT 1245.370 1320.745 1249.130 1321.025 ;
        RECT 1249.970 1320.745 1254.650 1321.025 ;
        RECT 1255.490 1320.745 1259.250 1321.025 ;
        RECT 1260.090 1320.745 1263.850 1321.025 ;
        RECT 1264.690 1320.745 1269.370 1321.025 ;
        RECT 1270.210 1320.745 1273.970 1321.025 ;
        RECT 1274.810 1320.745 1278.570 1321.025 ;
        RECT 1279.410 1320.745 1284.090 1321.025 ;
        RECT 1284.930 1320.745 1288.690 1321.025 ;
        RECT 1289.530 1320.745 1294.210 1321.025 ;
        RECT 1295.050 1320.745 1298.810 1321.025 ;
        RECT 1299.650 1320.745 1303.410 1321.025 ;
        RECT 1304.250 1320.745 1308.930 1321.025 ;
        RECT 1309.770 1320.745 1313.530 1321.025 ;
        RECT 1314.370 1320.745 1318.130 1321.025 ;
        RECT 1318.970 1320.745 1323.650 1321.025 ;
        RECT 1324.490 1320.745 1328.250 1321.025 ;
        RECT 1329.090 1320.745 1333.770 1321.025 ;
        RECT 1334.610 1320.745 1338.370 1321.025 ;
        RECT 1339.210 1320.745 1342.970 1321.025 ;
        RECT 1343.810 1320.745 1348.490 1321.025 ;
        RECT 1349.330 1320.745 1353.090 1321.025 ;
        RECT 1353.930 1320.745 1357.690 1321.025 ;
        RECT 1358.530 1320.745 1363.210 1321.025 ;
        RECT 1364.050 1320.745 1367.810 1321.025 ;
        RECT 1368.650 1320.745 1373.330 1321.025 ;
        RECT 1374.170 1320.745 1377.930 1321.025 ;
        RECT 1378.770 1320.745 1382.530 1321.025 ;
        RECT 1383.370 1320.745 1388.050 1321.025 ;
        RECT 1388.890 1320.745 1392.650 1321.025 ;
        RECT 1393.490 1320.745 1397.250 1321.025 ;
        RECT 1398.090 1320.745 1402.770 1321.025 ;
        RECT 312.860 220.280 1403.320 1320.745 ;
        RECT 313.410 220.000 317.170 220.280 ;
        RECT 318.010 220.000 321.770 220.280 ;
        RECT 322.610 220.000 327.290 220.280 ;
        RECT 328.130 220.000 331.890 220.280 ;
        RECT 332.730 220.000 336.490 220.280 ;
        RECT 337.330 220.000 342.010 220.280 ;
        RECT 342.850 220.000 346.610 220.280 ;
        RECT 347.450 220.000 352.130 220.280 ;
        RECT 352.970 220.000 356.730 220.280 ;
        RECT 357.570 220.000 361.330 220.280 ;
        RECT 362.170 220.000 366.850 220.280 ;
        RECT 367.690 220.000 371.450 220.280 ;
        RECT 372.290 220.000 376.050 220.280 ;
        RECT 376.890 220.000 381.570 220.280 ;
        RECT 382.410 220.000 386.170 220.280 ;
        RECT 387.010 220.000 391.690 220.280 ;
        RECT 392.530 220.000 396.290 220.280 ;
        RECT 397.130 220.000 400.890 220.280 ;
        RECT 401.730 220.000 406.410 220.280 ;
        RECT 407.250 220.000 411.010 220.280 ;
        RECT 411.850 220.000 415.610 220.280 ;
        RECT 416.450 220.000 421.130 220.280 ;
        RECT 421.970 220.000 425.730 220.280 ;
        RECT 426.570 220.000 431.250 220.280 ;
        RECT 432.090 220.000 435.850 220.280 ;
        RECT 436.690 220.000 440.450 220.280 ;
        RECT 441.290 220.000 445.970 220.280 ;
        RECT 446.810 220.000 450.570 220.280 ;
        RECT 451.410 220.000 455.170 220.280 ;
        RECT 456.010 220.000 460.690 220.280 ;
        RECT 461.530 220.000 465.290 220.280 ;
        RECT 466.130 220.000 470.810 220.280 ;
        RECT 471.650 220.000 475.410 220.280 ;
        RECT 476.250 220.000 480.010 220.280 ;
        RECT 480.850 220.000 485.530 220.280 ;
        RECT 486.370 220.000 490.130 220.280 ;
        RECT 490.970 220.000 494.730 220.280 ;
        RECT 495.570 220.000 500.250 220.280 ;
        RECT 501.090 220.000 504.850 220.280 ;
        RECT 505.690 220.000 510.370 220.280 ;
        RECT 511.210 220.000 514.970 220.280 ;
        RECT 515.810 220.000 519.570 220.280 ;
        RECT 520.410 220.000 525.090 220.280 ;
        RECT 525.930 220.000 529.690 220.280 ;
        RECT 530.530 220.000 534.290 220.280 ;
        RECT 535.130 220.000 539.810 220.280 ;
        RECT 540.650 220.000 544.410 220.280 ;
        RECT 545.250 220.000 549.930 220.280 ;
        RECT 550.770 220.000 554.530 220.280 ;
        RECT 555.370 220.000 559.130 220.280 ;
        RECT 559.970 220.000 564.650 220.280 ;
        RECT 565.490 220.000 569.250 220.280 ;
        RECT 570.090 220.000 573.850 220.280 ;
        RECT 574.690 220.000 579.370 220.280 ;
        RECT 580.210 220.000 583.970 220.280 ;
        RECT 584.810 220.000 589.490 220.280 ;
        RECT 590.330 220.000 594.090 220.280 ;
        RECT 594.930 220.000 598.690 220.280 ;
        RECT 599.530 220.000 604.210 220.280 ;
        RECT 605.050 220.000 608.810 220.280 ;
        RECT 609.650 220.000 613.410 220.280 ;
        RECT 614.250 220.000 618.930 220.280 ;
        RECT 619.770 220.000 623.530 220.280 ;
        RECT 624.370 220.000 629.050 220.280 ;
        RECT 629.890 220.000 633.650 220.280 ;
        RECT 634.490 220.000 638.250 220.280 ;
        RECT 639.090 220.000 643.770 220.280 ;
        RECT 644.610 220.000 648.370 220.280 ;
        RECT 649.210 220.000 652.970 220.280 ;
        RECT 653.810 220.000 658.490 220.280 ;
        RECT 659.330 220.000 663.090 220.280 ;
        RECT 663.930 220.000 668.610 220.280 ;
        RECT 669.450 220.000 673.210 220.280 ;
        RECT 674.050 220.000 677.810 220.280 ;
        RECT 678.650 220.000 683.330 220.280 ;
        RECT 684.170 220.000 687.930 220.280 ;
        RECT 688.770 220.000 692.530 220.280 ;
        RECT 693.370 220.000 698.050 220.280 ;
        RECT 698.890 220.000 702.650 220.280 ;
        RECT 703.490 220.000 708.170 220.280 ;
        RECT 709.010 220.000 712.770 220.280 ;
        RECT 713.610 220.000 717.370 220.280 ;
        RECT 718.210 220.000 722.890 220.280 ;
        RECT 723.730 220.000 727.490 220.280 ;
        RECT 728.330 220.000 732.090 220.280 ;
        RECT 732.930 220.000 737.610 220.280 ;
        RECT 738.450 220.000 742.210 220.280 ;
        RECT 743.050 220.000 747.730 220.280 ;
        RECT 748.570 220.000 752.330 220.280 ;
        RECT 753.170 220.000 756.930 220.280 ;
        RECT 757.770 220.000 762.450 220.280 ;
        RECT 763.290 220.000 767.050 220.280 ;
        RECT 767.890 220.000 771.650 220.280 ;
        RECT 772.490 220.000 777.170 220.280 ;
        RECT 778.010 220.000 781.770 220.280 ;
        RECT 782.610 220.000 787.290 220.280 ;
        RECT 788.130 220.000 791.890 220.280 ;
        RECT 792.730 220.000 796.490 220.280 ;
        RECT 797.330 220.000 802.010 220.280 ;
        RECT 802.850 220.000 806.610 220.280 ;
        RECT 807.450 220.000 811.210 220.280 ;
        RECT 812.050 220.000 816.730 220.280 ;
        RECT 817.570 220.000 821.330 220.280 ;
        RECT 822.170 220.000 826.850 220.280 ;
        RECT 827.690 220.000 831.450 220.280 ;
        RECT 832.290 220.000 836.050 220.280 ;
        RECT 836.890 220.000 841.570 220.280 ;
        RECT 842.410 220.000 846.170 220.280 ;
        RECT 847.010 220.000 850.770 220.280 ;
        RECT 851.610 220.000 856.290 220.280 ;
        RECT 857.130 220.000 860.890 220.280 ;
        RECT 861.730 220.000 866.410 220.280 ;
        RECT 867.250 220.000 871.010 220.280 ;
        RECT 871.850 220.000 875.610 220.280 ;
        RECT 876.450 220.000 881.130 220.280 ;
        RECT 881.970 220.000 885.730 220.280 ;
        RECT 886.570 220.000 890.330 220.280 ;
        RECT 891.170 220.000 895.850 220.280 ;
        RECT 896.690 220.000 900.450 220.280 ;
        RECT 901.290 220.000 905.970 220.280 ;
        RECT 906.810 220.000 910.570 220.280 ;
        RECT 911.410 220.000 915.170 220.280 ;
        RECT 916.010 220.000 920.690 220.280 ;
        RECT 921.530 220.000 925.290 220.280 ;
        RECT 926.130 220.000 929.890 220.280 ;
        RECT 930.730 220.000 935.410 220.280 ;
        RECT 936.250 220.000 940.010 220.280 ;
        RECT 940.850 220.000 945.530 220.280 ;
        RECT 946.370 220.000 950.130 220.280 ;
        RECT 950.970 220.000 954.730 220.280 ;
        RECT 955.570 220.000 960.250 220.280 ;
        RECT 961.090 220.000 964.850 220.280 ;
        RECT 965.690 220.000 969.450 220.280 ;
        RECT 970.290 220.000 974.970 220.280 ;
        RECT 975.810 220.000 979.570 220.280 ;
        RECT 980.410 220.000 985.090 220.280 ;
        RECT 985.930 220.000 989.690 220.280 ;
        RECT 990.530 220.000 994.290 220.280 ;
        RECT 995.130 220.000 999.810 220.280 ;
        RECT 1000.650 220.000 1004.410 220.280 ;
        RECT 1005.250 220.000 1009.010 220.280 ;
        RECT 1009.850 220.000 1014.530 220.280 ;
        RECT 1015.370 220.000 1019.130 220.280 ;
        RECT 1019.970 220.000 1024.650 220.280 ;
        RECT 1025.490 220.000 1029.250 220.280 ;
        RECT 1030.090 220.000 1033.850 220.280 ;
        RECT 1034.690 220.000 1039.370 220.280 ;
        RECT 1040.210 220.000 1043.970 220.280 ;
        RECT 1044.810 220.000 1048.570 220.280 ;
        RECT 1049.410 220.000 1054.090 220.280 ;
        RECT 1054.930 220.000 1058.690 220.280 ;
        RECT 1059.530 220.000 1064.210 220.280 ;
        RECT 1065.050 220.000 1068.810 220.280 ;
        RECT 1069.650 220.000 1073.410 220.280 ;
        RECT 1074.250 220.000 1078.930 220.280 ;
        RECT 1079.770 220.000 1083.530 220.280 ;
        RECT 1084.370 220.000 1088.130 220.280 ;
        RECT 1088.970 220.000 1093.650 220.280 ;
        RECT 1094.490 220.000 1098.250 220.280 ;
        RECT 1099.090 220.000 1103.770 220.280 ;
        RECT 1104.610 220.000 1108.370 220.280 ;
        RECT 1109.210 220.000 1112.970 220.280 ;
        RECT 1113.810 220.000 1118.490 220.280 ;
        RECT 1119.330 220.000 1123.090 220.280 ;
        RECT 1123.930 220.000 1127.690 220.280 ;
        RECT 1128.530 220.000 1133.210 220.280 ;
        RECT 1134.050 220.000 1137.810 220.280 ;
        RECT 1138.650 220.000 1143.330 220.280 ;
        RECT 1144.170 220.000 1147.930 220.280 ;
        RECT 1148.770 220.000 1152.530 220.280 ;
        RECT 1153.370 220.000 1158.050 220.280 ;
        RECT 1158.890 220.000 1162.650 220.280 ;
        RECT 1163.490 220.000 1167.250 220.280 ;
        RECT 1168.090 220.000 1172.770 220.280 ;
        RECT 1173.610 220.000 1177.370 220.280 ;
        RECT 1178.210 220.000 1182.890 220.280 ;
        RECT 1183.730 220.000 1187.490 220.280 ;
        RECT 1188.330 220.000 1192.090 220.280 ;
        RECT 1192.930 220.000 1197.610 220.280 ;
        RECT 1198.450 220.000 1202.210 220.280 ;
        RECT 1203.050 220.000 1206.810 220.280 ;
        RECT 1207.650 220.000 1212.330 220.280 ;
        RECT 1213.170 220.000 1216.930 220.280 ;
        RECT 1217.770 220.000 1222.450 220.280 ;
        RECT 1223.290 220.000 1227.050 220.280 ;
        RECT 1227.890 220.000 1231.650 220.280 ;
        RECT 1232.490 220.000 1237.170 220.280 ;
        RECT 1238.010 220.000 1241.770 220.280 ;
        RECT 1242.610 220.000 1246.370 220.280 ;
        RECT 1247.210 220.000 1251.890 220.280 ;
        RECT 1252.730 220.000 1256.490 220.280 ;
        RECT 1257.330 220.000 1262.010 220.280 ;
        RECT 1262.850 220.000 1266.610 220.280 ;
        RECT 1267.450 220.000 1271.210 220.280 ;
        RECT 1272.050 220.000 1276.730 220.280 ;
        RECT 1277.570 220.000 1281.330 220.280 ;
        RECT 1282.170 220.000 1285.930 220.280 ;
        RECT 1286.770 220.000 1291.450 220.280 ;
        RECT 1292.290 220.000 1296.050 220.280 ;
        RECT 1296.890 220.000 1301.570 220.280 ;
        RECT 1302.410 220.000 1306.170 220.280 ;
        RECT 1307.010 220.000 1310.770 220.280 ;
        RECT 1311.610 220.000 1316.290 220.280 ;
        RECT 1317.130 220.000 1320.890 220.280 ;
        RECT 1321.730 220.000 1325.490 220.280 ;
        RECT 1326.330 220.000 1331.010 220.280 ;
        RECT 1331.850 220.000 1335.610 220.280 ;
        RECT 1336.450 220.000 1341.130 220.280 ;
        RECT 1341.970 220.000 1345.730 220.280 ;
        RECT 1346.570 220.000 1350.330 220.280 ;
        RECT 1351.170 220.000 1355.850 220.280 ;
        RECT 1356.690 220.000 1360.450 220.280 ;
        RECT 1361.290 220.000 1365.050 220.280 ;
        RECT 1365.890 220.000 1370.570 220.280 ;
        RECT 1371.410 220.000 1375.170 220.280 ;
        RECT 1376.010 220.000 1380.690 220.280 ;
        RECT 1381.530 220.000 1385.290 220.280 ;
        RECT 1386.130 220.000 1389.890 220.280 ;
        RECT 1390.730 220.000 1395.410 220.280 ;
        RECT 1396.250 220.000 1400.010 220.280 ;
        RECT 1400.850 220.000 1403.320 220.280 ;
      LAYER met2 ;
        RECT 312.850 216.000 313.130 220.000 ;
        RECT 327.570 216.000 327.850 220.000 ;
        RECT 332.170 216.000 332.450 220.000 ;
        RECT 336.770 216.000 337.050 220.000 ;
        RECT 361.610 216.000 361.890 220.000 ;
        RECT 367.130 216.000 367.410 220.000 ;
        RECT 376.330 216.000 376.610 220.000 ;
        RECT 381.850 216.000 382.130 220.000 ;
        RECT 386.450 216.000 386.730 220.000 ;
        RECT 391.970 216.000 392.250 220.000 ;
        RECT 401.170 216.000 401.450 220.000 ;
        RECT 426.010 216.000 426.290 220.000 ;
        RECT 450.850 216.000 451.130 220.000 ;
        RECT 465.570 216.000 465.850 220.000 ;
        RECT 490.410 216.000 490.690 220.000 ;
        RECT 510.650 216.000 510.930 220.000 ;
        RECT 525.370 216.000 525.650 220.000 ;
        RECT 540.090 216.000 540.370 220.000 ;
        RECT 550.210 216.000 550.490 220.000 ;
        RECT 569.530 216.000 569.810 220.000 ;
        RECT 579.650 216.000 579.930 220.000 ;
        RECT 584.250 216.000 584.530 220.000 ;
        RECT 609.090 216.000 609.370 220.000 ;
        RECT 623.810 216.000 624.090 220.000 ;
        RECT 668.890 216.000 669.170 220.000 ;
        RECT 688.210 216.000 688.490 220.000 ;
        RECT 752.610 216.000 752.890 220.000 ;
        RECT 771.930 216.000 772.210 220.000 ;
        RECT 782.050 216.000 782.330 220.000 ;
        RECT 796.770 216.000 797.050 220.000 ;
        RECT 827.130 216.000 827.410 220.000 ;
        RECT 831.730 216.000 832.010 220.000 ;
        RECT 875.890 216.000 876.170 220.000 ;
        RECT 881.410 216.000 881.690 220.000 ;
        RECT 886.010 216.000 886.290 220.000 ;
        RECT 940.290 216.000 940.570 220.000 ;
        RECT 960.530 216.000 960.810 220.000 ;
        RECT 969.730 216.000 970.010 220.000 ;
        RECT 1004.690 216.000 1004.970 220.000 ;
        RECT 1009.290 216.000 1009.570 220.000 ;
        RECT 1034.130 216.000 1034.410 220.000 ;
        RECT 1044.250 216.000 1044.530 220.000 ;
        RECT 1088.410 216.000 1088.690 220.000 ;
        RECT 1093.930 216.000 1094.210 220.000 ;
        RECT 1113.250 216.000 1113.530 220.000 ;
        RECT 1133.490 216.000 1133.770 220.000 ;
        RECT 1138.090 216.000 1138.370 220.000 ;
        RECT 1143.610 216.000 1143.890 220.000 ;
        RECT 1158.330 216.000 1158.610 220.000 ;
        RECT 1162.930 216.000 1163.210 220.000 ;
        RECT 1183.170 216.000 1183.450 220.000 ;
        RECT 1296.330 216.000 1296.610 220.000 ;
        RECT 1301.850 216.000 1302.130 220.000 ;
        RECT 1311.050 216.000 1311.330 220.000 ;
        RECT 1316.570 216.000 1316.850 220.000 ;
        RECT 1360.730 216.000 1361.010 220.000 ;
        RECT 1365.330 216.000 1365.610 220.000 ;
        RECT 1375.450 216.000 1375.730 220.000 ;
        RECT 1385.570 216.000 1385.850 220.000 ;
        RECT 1400.290 216.000 1400.570 220.000 ;
      LAYER met3 ;
        RECT 310.000 1316.280 314.000 1316.880 ;
      LAYER met3 ;
        RECT 314.400 1315.880 1403.905 1316.745 ;
      LAYER met3 ;
        RECT 1404.305 1316.280 1408.305 1316.880 ;
      LAYER met3 ;
        RECT 313.990 1309.120 1404.305 1315.880 ;
      LAYER met3 ;
        RECT 310.000 1308.120 314.000 1308.720 ;
      LAYER met3 ;
        RECT 314.400 1307.720 1403.905 1309.120 ;
        RECT 313.990 1302.320 1404.305 1307.720 ;
        RECT 314.400 1300.920 1403.905 1302.320 ;
      LAYER met3 ;
        RECT 1404.305 1301.320 1408.305 1301.920 ;
      LAYER met3 ;
        RECT 313.990 1295.520 1404.305 1300.920 ;
      LAYER met3 ;
        RECT 310.000 1294.520 314.000 1295.120 ;
      LAYER met3 ;
        RECT 314.400 1294.120 1403.905 1295.520 ;
      LAYER met3 ;
        RECT 1404.305 1294.520 1408.305 1295.120 ;
      LAYER met3 ;
        RECT 313.990 1287.360 1404.305 1294.120 ;
        RECT 314.400 1285.960 1403.905 1287.360 ;
      LAYER met3 ;
        RECT 1404.305 1286.360 1408.305 1286.960 ;
      LAYER met3 ;
        RECT 313.990 1280.560 1404.305 1285.960 ;
      LAYER met3 ;
        RECT 310.000 1279.560 314.000 1280.160 ;
      LAYER met3 ;
        RECT 314.400 1279.160 1403.905 1280.560 ;
        RECT 313.990 1273.760 1404.305 1279.160 ;
      LAYER met3 ;
        RECT 310.000 1272.760 314.000 1273.360 ;
      LAYER met3 ;
        RECT 314.400 1272.360 1403.905 1273.760 ;
      LAYER met3 ;
        RECT 1404.305 1272.760 1408.305 1273.360 ;
      LAYER met3 ;
        RECT 313.990 1265.600 1404.305 1272.360 ;
        RECT 314.400 1264.200 1403.905 1265.600 ;
        RECT 313.990 1258.800 1404.305 1264.200 ;
        RECT 314.400 1257.400 1403.905 1258.800 ;
        RECT 313.990 1250.640 1404.305 1257.400 ;
        RECT 314.400 1249.240 1403.905 1250.640 ;
        RECT 313.990 1243.840 1404.305 1249.240 ;
        RECT 314.400 1242.440 1403.905 1243.840 ;
        RECT 313.990 1237.040 1404.305 1242.440 ;
        RECT 314.400 1235.640 1403.905 1237.040 ;
      LAYER met3 ;
        RECT 1404.305 1236.040 1408.305 1236.640 ;
      LAYER met3 ;
        RECT 313.990 1228.880 1404.305 1235.640 ;
      LAYER met3 ;
        RECT 310.000 1227.880 314.000 1228.480 ;
      LAYER met3 ;
        RECT 314.400 1227.480 1403.905 1228.880 ;
        RECT 313.990 1222.080 1404.305 1227.480 ;
        RECT 314.400 1220.680 1403.905 1222.080 ;
        RECT 313.990 1215.280 1404.305 1220.680 ;
      LAYER met3 ;
        RECT 310.000 1214.280 314.000 1214.880 ;
      LAYER met3 ;
        RECT 314.400 1213.880 1403.905 1215.280 ;
      LAYER met3 ;
        RECT 1404.305 1214.280 1408.305 1214.880 ;
      LAYER met3 ;
        RECT 313.990 1207.120 1404.305 1213.880 ;
      LAYER met3 ;
        RECT 310.000 1206.120 314.000 1206.720 ;
      LAYER met3 ;
        RECT 314.400 1205.720 1403.905 1207.120 ;
        RECT 313.990 1200.320 1404.305 1205.720 ;
        RECT 314.400 1198.920 1403.905 1200.320 ;
      LAYER met3 ;
        RECT 1404.305 1199.320 1408.305 1199.920 ;
      LAYER met3 ;
        RECT 313.990 1192.160 1404.305 1198.920 ;
        RECT 314.400 1190.760 1403.905 1192.160 ;
        RECT 313.990 1185.360 1404.305 1190.760 ;
        RECT 314.400 1183.960 1403.905 1185.360 ;
      LAYER met3 ;
        RECT 1404.305 1184.360 1408.305 1184.960 ;
      LAYER met3 ;
        RECT 313.990 1178.560 1404.305 1183.960 ;
      LAYER met3 ;
        RECT 310.000 1177.560 314.000 1178.160 ;
      LAYER met3 ;
        RECT 314.400 1177.160 1403.905 1178.560 ;
        RECT 313.990 1170.400 1404.305 1177.160 ;
        RECT 314.400 1169.000 1403.905 1170.400 ;
        RECT 313.990 1163.600 1404.305 1169.000 ;
      LAYER met3 ;
        RECT 310.000 1162.600 314.000 1163.200 ;
      LAYER met3 ;
        RECT 314.400 1162.200 1403.905 1163.600 ;
      LAYER met3 ;
        RECT 1404.305 1162.600 1408.305 1163.200 ;
      LAYER met3 ;
        RECT 313.990 1156.800 1404.305 1162.200 ;
      LAYER met3 ;
        RECT 310.000 1155.800 314.000 1156.400 ;
      LAYER met3 ;
        RECT 314.400 1155.400 1403.905 1156.800 ;
      LAYER met3 ;
        RECT 1404.305 1155.800 1408.305 1156.400 ;
      LAYER met3 ;
        RECT 313.990 1148.640 1404.305 1155.400 ;
        RECT 314.400 1147.240 1403.905 1148.640 ;
      LAYER met3 ;
        RECT 1404.305 1147.640 1408.305 1148.240 ;
      LAYER met3 ;
        RECT 313.990 1141.840 1404.305 1147.240 ;
        RECT 314.400 1140.440 1403.905 1141.840 ;
        RECT 313.990 1133.680 1404.305 1140.440 ;
      LAYER met3 ;
        RECT 310.000 1132.680 314.000 1133.280 ;
      LAYER met3 ;
        RECT 314.400 1132.280 1403.905 1133.680 ;
        RECT 313.990 1126.880 1404.305 1132.280 ;
      LAYER met3 ;
        RECT 310.000 1125.880 314.000 1126.480 ;
      LAYER met3 ;
        RECT 314.400 1125.480 1403.905 1126.880 ;
        RECT 313.990 1120.080 1404.305 1125.480 ;
        RECT 314.400 1118.680 1403.905 1120.080 ;
      LAYER met3 ;
        RECT 1404.305 1119.080 1408.305 1119.680 ;
      LAYER met3 ;
        RECT 313.990 1111.920 1404.305 1118.680 ;
        RECT 314.400 1110.520 1403.905 1111.920 ;
      LAYER met3 ;
        RECT 1404.305 1110.920 1408.305 1111.520 ;
      LAYER met3 ;
        RECT 313.990 1105.120 1404.305 1110.520 ;
        RECT 314.400 1103.720 1403.905 1105.120 ;
      LAYER met3 ;
        RECT 1404.305 1104.120 1408.305 1104.720 ;
      LAYER met3 ;
        RECT 313.990 1098.320 1404.305 1103.720 ;
        RECT 314.400 1096.920 1403.905 1098.320 ;
        RECT 313.990 1090.160 1404.305 1096.920 ;
        RECT 314.400 1088.760 1403.905 1090.160 ;
        RECT 313.990 1083.360 1404.305 1088.760 ;
        RECT 314.400 1081.960 1403.905 1083.360 ;
        RECT 313.990 1075.200 1404.305 1081.960 ;
        RECT 314.400 1073.800 1403.905 1075.200 ;
        RECT 313.990 1068.400 1404.305 1073.800 ;
        RECT 314.400 1067.000 1403.905 1068.400 ;
        RECT 313.990 1061.600 1404.305 1067.000 ;
        RECT 314.400 1060.200 1403.905 1061.600 ;
        RECT 313.990 1053.440 1404.305 1060.200 ;
        RECT 314.400 1052.040 1403.905 1053.440 ;
      LAYER met3 ;
        RECT 1404.305 1052.440 1408.305 1053.040 ;
      LAYER met3 ;
        RECT 313.990 1046.640 1404.305 1052.040 ;
      LAYER met3 ;
        RECT 310.000 1045.640 314.000 1046.240 ;
      LAYER met3 ;
        RECT 314.400 1045.240 1403.905 1046.640 ;
        RECT 313.990 1039.840 1404.305 1045.240 ;
      LAYER met3 ;
        RECT 310.000 1038.840 314.000 1039.440 ;
      LAYER met3 ;
        RECT 314.400 1038.440 1403.905 1039.840 ;
        RECT 313.990 1031.680 1404.305 1038.440 ;
        RECT 314.400 1030.280 1403.905 1031.680 ;
      LAYER met3 ;
        RECT 1404.305 1030.680 1408.305 1031.280 ;
      LAYER met3 ;
        RECT 313.990 1024.880 1404.305 1030.280 ;
      LAYER met3 ;
        RECT 310.000 1023.880 314.000 1024.480 ;
      LAYER met3 ;
        RECT 314.400 1023.480 1403.905 1024.880 ;
        RECT 313.990 1016.720 1404.305 1023.480 ;
        RECT 314.400 1015.320 1403.905 1016.720 ;
      LAYER met3 ;
        RECT 1404.305 1015.720 1408.305 1016.320 ;
      LAYER met3 ;
        RECT 313.990 1009.920 1404.305 1015.320 ;
      LAYER met3 ;
        RECT 310.000 1008.920 314.000 1009.520 ;
      LAYER met3 ;
        RECT 314.400 1008.520 1403.905 1009.920 ;
        RECT 313.990 1003.120 1404.305 1008.520 ;
        RECT 314.400 1001.720 1403.905 1003.120 ;
      LAYER met3 ;
        RECT 1404.305 1002.120 1408.305 1002.720 ;
      LAYER met3 ;
        RECT 313.990 994.960 1404.305 1001.720 ;
        RECT 314.400 993.560 1403.905 994.960 ;
        RECT 313.990 988.160 1404.305 993.560 ;
      LAYER met3 ;
        RECT 310.000 987.160 314.000 987.760 ;
      LAYER met3 ;
        RECT 314.400 986.760 1403.905 988.160 ;
        RECT 313.990 981.360 1404.305 986.760 ;
      LAYER met3 ;
        RECT 310.000 980.360 314.000 980.960 ;
      LAYER met3 ;
        RECT 314.400 979.960 1403.905 981.360 ;
      LAYER met3 ;
        RECT 1404.305 980.360 1408.305 980.960 ;
      LAYER met3 ;
        RECT 313.990 973.200 1404.305 979.960 ;
        RECT 314.400 971.800 1403.905 973.200 ;
        RECT 313.990 966.400 1404.305 971.800 ;
        RECT 314.400 965.000 1403.905 966.400 ;
        RECT 313.990 958.240 1404.305 965.000 ;
        RECT 314.400 956.840 1403.905 958.240 ;
        RECT 313.990 951.440 1404.305 956.840 ;
        RECT 314.400 950.040 1403.905 951.440 ;
        RECT 313.990 944.640 1404.305 950.040 ;
        RECT 314.400 943.240 1403.905 944.640 ;
        RECT 313.990 936.480 1404.305 943.240 ;
        RECT 314.400 935.080 1403.905 936.480 ;
      LAYER met3 ;
        RECT 1404.305 935.480 1408.305 936.080 ;
      LAYER met3 ;
        RECT 313.990 929.680 1404.305 935.080 ;
        RECT 314.400 928.280 1403.905 929.680 ;
        RECT 313.990 922.880 1404.305 928.280 ;
      LAYER met3 ;
        RECT 310.000 921.880 314.000 922.480 ;
      LAYER met3 ;
        RECT 314.400 921.480 1403.905 922.880 ;
        RECT 313.990 914.720 1404.305 921.480 ;
        RECT 314.400 913.320 1403.905 914.720 ;
        RECT 313.990 907.920 1404.305 913.320 ;
        RECT 314.400 906.520 1403.905 907.920 ;
      LAYER met3 ;
        RECT 1404.305 906.920 1408.305 907.520 ;
      LAYER met3 ;
        RECT 313.990 899.760 1404.305 906.520 ;
      LAYER met3 ;
        RECT 310.000 898.760 314.000 899.360 ;
      LAYER met3 ;
        RECT 314.400 898.360 1403.905 899.760 ;
        RECT 313.990 892.960 1404.305 898.360 ;
      LAYER met3 ;
        RECT 310.000 891.960 314.000 892.560 ;
      LAYER met3 ;
        RECT 314.400 891.560 1403.905 892.960 ;
      LAYER met3 ;
        RECT 1404.305 891.960 1408.305 892.560 ;
      LAYER met3 ;
        RECT 313.990 886.160 1404.305 891.560 ;
      LAYER met3 ;
        RECT 310.000 885.160 314.000 885.760 ;
      LAYER met3 ;
        RECT 314.400 884.760 1403.905 886.160 ;
        RECT 313.990 878.000 1404.305 884.760 ;
        RECT 314.400 876.600 1403.905 878.000 ;
      LAYER met3 ;
        RECT 1404.305 877.000 1408.305 877.600 ;
      LAYER met3 ;
        RECT 313.990 871.200 1404.305 876.600 ;
        RECT 314.400 869.800 1403.905 871.200 ;
        RECT 313.990 864.400 1404.305 869.800 ;
        RECT 314.400 863.000 1403.905 864.400 ;
        RECT 313.990 856.240 1404.305 863.000 ;
        RECT 314.400 854.840 1403.905 856.240 ;
        RECT 313.990 849.440 1404.305 854.840 ;
      LAYER met3 ;
        RECT 310.000 848.440 314.000 849.040 ;
      LAYER met3 ;
        RECT 314.400 848.040 1403.905 849.440 ;
      LAYER met3 ;
        RECT 1404.305 848.440 1408.305 849.040 ;
      LAYER met3 ;
        RECT 313.990 841.280 1404.305 848.040 ;
        RECT 314.400 839.880 1403.905 841.280 ;
        RECT 313.990 834.480 1404.305 839.880 ;
      LAYER met3 ;
        RECT 310.000 833.480 314.000 834.080 ;
      LAYER met3 ;
        RECT 314.400 833.080 1403.905 834.480 ;
      LAYER met3 ;
        RECT 1404.305 833.480 1408.305 834.080 ;
      LAYER met3 ;
        RECT 313.990 827.680 1404.305 833.080 ;
        RECT 314.400 826.280 1403.905 827.680 ;
        RECT 313.990 819.520 1404.305 826.280 ;
        RECT 314.400 818.120 1403.905 819.520 ;
        RECT 313.990 812.720 1404.305 818.120 ;
      LAYER met3 ;
        RECT 310.000 811.720 314.000 812.320 ;
      LAYER met3 ;
        RECT 314.400 811.320 1403.905 812.720 ;
        RECT 313.990 805.920 1404.305 811.320 ;
        RECT 314.400 804.520 1403.905 805.920 ;
        RECT 313.990 797.760 1404.305 804.520 ;
        RECT 314.400 796.360 1403.905 797.760 ;
      LAYER met3 ;
        RECT 1404.305 796.760 1408.305 797.360 ;
      LAYER met3 ;
        RECT 313.990 790.960 1404.305 796.360 ;
        RECT 314.400 789.560 1403.905 790.960 ;
      LAYER met3 ;
        RECT 1404.305 789.960 1408.305 790.560 ;
      LAYER met3 ;
        RECT 313.990 782.800 1404.305 789.560 ;
      LAYER met3 ;
        RECT 310.000 781.800 314.000 782.400 ;
      LAYER met3 ;
        RECT 314.400 781.400 1403.905 782.800 ;
        RECT 313.990 776.000 1404.305 781.400 ;
      LAYER met3 ;
        RECT 310.000 775.000 314.000 775.600 ;
      LAYER met3 ;
        RECT 314.400 774.600 1403.905 776.000 ;
      LAYER met3 ;
        RECT 1404.305 775.000 1408.305 775.600 ;
      LAYER met3 ;
        RECT 313.990 769.200 1404.305 774.600 ;
        RECT 314.400 767.800 1403.905 769.200 ;
        RECT 313.990 761.040 1404.305 767.800 ;
      LAYER met3 ;
        RECT 310.000 760.040 314.000 760.640 ;
      LAYER met3 ;
        RECT 314.400 759.640 1403.905 761.040 ;
        RECT 313.990 754.240 1404.305 759.640 ;
        RECT 314.400 752.840 1403.905 754.240 ;
      LAYER met3 ;
        RECT 1404.305 753.240 1408.305 753.840 ;
      LAYER met3 ;
        RECT 313.990 747.440 1404.305 752.840 ;
        RECT 314.400 746.040 1403.905 747.440 ;
        RECT 313.990 739.280 1404.305 746.040 ;
        RECT 314.400 737.880 1403.905 739.280 ;
      LAYER met3 ;
        RECT 1404.305 738.280 1408.305 738.880 ;
      LAYER met3 ;
        RECT 313.990 732.480 1404.305 737.880 ;
        RECT 314.400 731.080 1403.905 732.480 ;
      LAYER met3 ;
        RECT 1404.305 731.480 1408.305 732.080 ;
      LAYER met3 ;
        RECT 313.990 724.320 1404.305 731.080 ;
        RECT 314.400 722.920 1403.905 724.320 ;
        RECT 313.990 717.520 1404.305 722.920 ;
        RECT 314.400 716.120 1403.905 717.520 ;
        RECT 313.990 710.720 1404.305 716.120 ;
        RECT 314.400 709.320 1403.905 710.720 ;
        RECT 313.990 702.560 1404.305 709.320 ;
      LAYER met3 ;
        RECT 310.000 701.560 314.000 702.160 ;
      LAYER met3 ;
        RECT 314.400 701.160 1403.905 702.560 ;
      LAYER met3 ;
        RECT 1404.305 701.560 1408.305 702.160 ;
      LAYER met3 ;
        RECT 313.990 695.760 1404.305 701.160 ;
      LAYER met3 ;
        RECT 310.000 694.760 314.000 695.360 ;
      LAYER met3 ;
        RECT 314.400 694.360 1403.905 695.760 ;
        RECT 313.990 688.960 1404.305 694.360 ;
        RECT 314.400 687.560 1403.905 688.960 ;
        RECT 313.990 680.800 1404.305 687.560 ;
      LAYER met3 ;
        RECT 310.000 679.800 314.000 680.400 ;
      LAYER met3 ;
        RECT 314.400 679.400 1403.905 680.800 ;
        RECT 313.990 674.000 1404.305 679.400 ;
      LAYER met3 ;
        RECT 310.000 673.000 314.000 673.600 ;
      LAYER met3 ;
        RECT 314.400 672.600 1403.905 674.000 ;
      LAYER met3 ;
        RECT 1404.305 673.000 1408.305 673.600 ;
      LAYER met3 ;
        RECT 313.990 665.840 1404.305 672.600 ;
        RECT 314.400 664.440 1403.905 665.840 ;
      LAYER met3 ;
        RECT 1404.305 664.840 1408.305 665.440 ;
      LAYER met3 ;
        RECT 313.990 659.040 1404.305 664.440 ;
        RECT 314.400 657.640 1403.905 659.040 ;
      LAYER met3 ;
        RECT 1404.305 658.040 1408.305 658.640 ;
      LAYER met3 ;
        RECT 313.990 652.240 1404.305 657.640 ;
        RECT 314.400 650.840 1403.905 652.240 ;
      LAYER met3 ;
        RECT 1404.305 651.240 1408.305 651.840 ;
      LAYER met3 ;
        RECT 313.990 644.080 1404.305 650.840 ;
        RECT 314.400 642.680 1403.905 644.080 ;
        RECT 313.990 637.280 1404.305 642.680 ;
      LAYER met3 ;
        RECT 310.000 636.280 314.000 636.880 ;
      LAYER met3 ;
        RECT 314.400 635.880 1403.905 637.280 ;
        RECT 313.990 630.480 1404.305 635.880 ;
      LAYER met3 ;
        RECT 310.000 629.480 314.000 630.080 ;
      LAYER met3 ;
        RECT 314.400 629.080 1403.905 630.480 ;
        RECT 313.990 622.320 1404.305 629.080 ;
      LAYER met3 ;
        RECT 310.000 621.320 314.000 621.920 ;
      LAYER met3 ;
        RECT 314.400 620.920 1403.905 622.320 ;
        RECT 313.990 615.520 1404.305 620.920 ;
        RECT 314.400 614.120 1403.905 615.520 ;
      LAYER met3 ;
        RECT 1404.305 614.520 1408.305 615.120 ;
      LAYER met3 ;
        RECT 313.990 607.360 1404.305 614.120 ;
        RECT 314.400 605.960 1403.905 607.360 ;
        RECT 313.990 600.560 1404.305 605.960 ;
        RECT 314.400 599.160 1403.905 600.560 ;
      LAYER met3 ;
        RECT 1404.305 599.560 1408.305 600.160 ;
      LAYER met3 ;
        RECT 313.990 593.760 1404.305 599.160 ;
        RECT 314.400 592.360 1403.905 593.760 ;
        RECT 313.990 585.600 1404.305 592.360 ;
      LAYER met3 ;
        RECT 310.000 584.600 314.000 585.200 ;
      LAYER met3 ;
        RECT 314.400 584.200 1403.905 585.600 ;
        RECT 313.990 578.800 1404.305 584.200 ;
      LAYER met3 ;
        RECT 310.000 577.800 314.000 578.400 ;
      LAYER met3 ;
        RECT 314.400 577.400 1403.905 578.800 ;
      LAYER met3 ;
        RECT 1404.305 577.800 1408.305 578.400 ;
      LAYER met3 ;
        RECT 313.990 572.000 1404.305 577.400 ;
      LAYER met3 ;
        RECT 310.000 571.000 314.000 571.600 ;
      LAYER met3 ;
        RECT 314.400 570.600 1403.905 572.000 ;
      LAYER met3 ;
        RECT 1404.305 571.000 1408.305 571.600 ;
      LAYER met3 ;
        RECT 313.990 563.840 1404.305 570.600 ;
        RECT 314.400 562.440 1403.905 563.840 ;
        RECT 313.990 557.040 1404.305 562.440 ;
        RECT 314.400 555.640 1403.905 557.040 ;
      LAYER met3 ;
        RECT 1404.305 556.040 1408.305 556.640 ;
      LAYER met3 ;
        RECT 313.990 548.880 1404.305 555.640 ;
        RECT 314.400 547.480 1403.905 548.880 ;
        RECT 313.990 542.080 1404.305 547.480 ;
      LAYER met3 ;
        RECT 310.000 541.080 314.000 541.680 ;
      LAYER met3 ;
        RECT 314.400 540.680 1403.905 542.080 ;
        RECT 313.990 535.280 1404.305 540.680 ;
        RECT 314.400 533.880 1403.905 535.280 ;
        RECT 313.990 527.120 1404.305 533.880 ;
        RECT 314.400 525.720 1403.905 527.120 ;
        RECT 313.990 520.320 1404.305 525.720 ;
        RECT 314.400 518.920 1403.905 520.320 ;
        RECT 313.990 513.520 1404.305 518.920 ;
      LAYER met3 ;
        RECT 310.000 512.520 314.000 513.120 ;
      LAYER met3 ;
        RECT 314.400 512.120 1403.905 513.520 ;
      LAYER met3 ;
        RECT 1404.305 512.520 1408.305 513.120 ;
      LAYER met3 ;
        RECT 313.990 505.360 1404.305 512.120 ;
        RECT 314.400 503.960 1403.905 505.360 ;
        RECT 313.990 498.560 1404.305 503.960 ;
      LAYER met3 ;
        RECT 310.000 497.560 314.000 498.160 ;
      LAYER met3 ;
        RECT 314.400 497.160 1403.905 498.560 ;
        RECT 313.990 490.400 1404.305 497.160 ;
        RECT 314.400 489.000 1403.905 490.400 ;
        RECT 313.990 483.600 1404.305 489.000 ;
      LAYER met3 ;
        RECT 310.000 482.600 314.000 483.200 ;
      LAYER met3 ;
        RECT 314.400 482.200 1403.905 483.600 ;
        RECT 313.990 476.800 1404.305 482.200 ;
        RECT 314.400 475.400 1403.905 476.800 ;
        RECT 313.990 468.640 1404.305 475.400 ;
      LAYER met3 ;
        RECT 310.000 467.640 314.000 468.240 ;
      LAYER met3 ;
        RECT 314.400 467.240 1403.905 468.640 ;
        RECT 313.990 461.840 1404.305 467.240 ;
      LAYER met3 ;
        RECT 310.000 460.840 314.000 461.440 ;
      LAYER met3 ;
        RECT 314.400 460.440 1403.905 461.840 ;
        RECT 313.990 455.040 1404.305 460.440 ;
        RECT 314.400 453.640 1403.905 455.040 ;
        RECT 313.990 446.880 1404.305 453.640 ;
      LAYER met3 ;
        RECT 310.000 445.880 314.000 446.480 ;
      LAYER met3 ;
        RECT 314.400 445.480 1403.905 446.880 ;
        RECT 313.990 440.080 1404.305 445.480 ;
        RECT 314.400 438.680 1403.905 440.080 ;
        RECT 313.990 431.920 1404.305 438.680 ;
        RECT 314.400 430.520 1403.905 431.920 ;
        RECT 313.990 425.120 1404.305 430.520 ;
      LAYER met3 ;
        RECT 310.000 424.120 314.000 424.720 ;
      LAYER met3 ;
        RECT 314.400 423.720 1403.905 425.120 ;
        RECT 313.990 418.320 1404.305 423.720 ;
        RECT 314.400 416.920 1403.905 418.320 ;
        RECT 313.990 410.160 1404.305 416.920 ;
        RECT 314.400 408.760 1403.905 410.160 ;
        RECT 313.990 403.360 1404.305 408.760 ;
        RECT 314.400 401.960 1403.905 403.360 ;
        RECT 313.990 396.560 1404.305 401.960 ;
        RECT 314.400 395.200 1404.305 396.560 ;
        RECT 314.400 395.160 1403.905 395.200 ;
        RECT 313.990 393.800 1403.905 395.160 ;
        RECT 313.990 388.400 1404.305 393.800 ;
        RECT 314.400 387.000 1403.905 388.400 ;
      LAYER met3 ;
        RECT 1404.305 387.400 1408.305 388.000 ;
      LAYER met3 ;
        RECT 313.990 381.600 1404.305 387.000 ;
        RECT 314.400 380.200 1403.905 381.600 ;
        RECT 313.990 373.440 1404.305 380.200 ;
        RECT 314.400 372.040 1403.905 373.440 ;
        RECT 313.990 366.640 1404.305 372.040 ;
      LAYER met3 ;
        RECT 310.000 365.640 314.000 366.240 ;
      LAYER met3 ;
        RECT 314.400 365.240 1403.905 366.640 ;
      LAYER met3 ;
        RECT 1404.305 365.640 1408.305 366.240 ;
      LAYER met3 ;
        RECT 313.990 359.840 1404.305 365.240 ;
      LAYER met3 ;
        RECT 310.000 358.840 314.000 359.440 ;
      LAYER met3 ;
        RECT 314.400 358.440 1403.905 359.840 ;
        RECT 313.990 351.680 1404.305 358.440 ;
        RECT 314.400 350.280 1403.905 351.680 ;
      LAYER met3 ;
        RECT 1404.305 350.680 1408.305 351.280 ;
      LAYER met3 ;
        RECT 313.990 344.880 1404.305 350.280 ;
      LAYER met3 ;
        RECT 310.000 343.880 314.000 344.480 ;
      LAYER met3 ;
        RECT 314.400 343.480 1403.905 344.880 ;
        RECT 313.990 338.080 1404.305 343.480 ;
      LAYER met3 ;
        RECT 310.000 337.080 314.000 337.680 ;
      LAYER met3 ;
        RECT 314.400 336.720 1404.305 338.080 ;
        RECT 314.400 336.680 1403.905 336.720 ;
        RECT 313.990 335.320 1403.905 336.680 ;
      LAYER met3 ;
        RECT 1404.305 335.720 1408.305 336.320 ;
      LAYER met3 ;
        RECT 313.990 329.920 1404.305 335.320 ;
        RECT 314.400 328.520 1403.905 329.920 ;
        RECT 313.990 323.120 1404.305 328.520 ;
        RECT 314.400 321.720 1403.905 323.120 ;
        RECT 313.990 314.960 1404.305 321.720 ;
      LAYER met3 ;
        RECT 310.000 313.960 314.000 314.560 ;
      LAYER met3 ;
        RECT 314.400 313.560 1403.905 314.960 ;
        RECT 313.990 308.160 1404.305 313.560 ;
        RECT 314.400 306.760 1403.905 308.160 ;
        RECT 313.990 301.360 1404.305 306.760 ;
        RECT 314.400 299.960 1403.905 301.360 ;
        RECT 313.990 293.200 1404.305 299.960 ;
        RECT 314.400 291.800 1403.905 293.200 ;
        RECT 313.990 286.400 1404.305 291.800 ;
      LAYER met3 ;
        RECT 310.000 285.400 314.000 286.000 ;
      LAYER met3 ;
        RECT 314.400 285.000 1403.905 286.400 ;
      LAYER met3 ;
        RECT 1404.305 285.400 1408.305 286.000 ;
      LAYER met3 ;
        RECT 313.990 279.600 1404.305 285.000 ;
      LAYER met3 ;
        RECT 310.000 278.600 314.000 279.200 ;
      LAYER met3 ;
        RECT 314.400 278.240 1404.305 279.600 ;
        RECT 314.400 278.200 1403.905 278.240 ;
        RECT 313.990 276.840 1403.905 278.200 ;
      LAYER met3 ;
        RECT 1404.305 277.240 1408.305 277.840 ;
      LAYER met3 ;
        RECT 313.990 271.440 1404.305 276.840 ;
        RECT 314.400 270.040 1403.905 271.440 ;
      LAYER met3 ;
        RECT 1404.305 270.440 1408.305 271.040 ;
      LAYER met3 ;
        RECT 313.990 264.640 1404.305 270.040 ;
      LAYER met3 ;
        RECT 310.000 263.640 314.000 264.240 ;
      LAYER met3 ;
        RECT 314.400 263.240 1403.905 264.640 ;
        RECT 313.990 256.480 1404.305 263.240 ;
      LAYER met3 ;
        RECT 310.000 255.480 314.000 256.080 ;
      LAYER met3 ;
        RECT 314.400 255.080 1403.905 256.480 ;
        RECT 313.990 249.680 1404.305 255.080 ;
        RECT 314.400 248.280 1403.905 249.680 ;
      LAYER met3 ;
        RECT 1404.305 248.680 1408.305 249.280 ;
      LAYER met3 ;
        RECT 313.990 242.880 1404.305 248.280 ;
        RECT 314.400 241.480 1403.905 242.880 ;
      LAYER met3 ;
        RECT 1404.305 241.880 1408.305 242.480 ;
      LAYER met3 ;
        RECT 313.990 234.720 1404.305 241.480 ;
        RECT 314.400 233.320 1403.905 234.720 ;
        RECT 313.990 227.920 1404.305 233.320 ;
        RECT 314.400 226.520 1403.905 227.920 ;
        RECT 313.990 220.255 1404.305 226.520 ;
      LAYER met4 ;
        RECT 325.015 226.640 1392.545 1312.400 ;
      LAYER met5 ;
        RECT 315.520 1182.380 1402.500 1239.760 ;
        RECT 315.520 1092.380 1402.500 1179.380 ;
        RECT 315.520 1002.380 1402.500 1089.380 ;
        RECT 315.520 912.380 1402.500 999.380 ;
        RECT 315.520 822.380 1402.500 909.380 ;
        RECT 315.520 732.380 1402.500 819.380 ;
        RECT 315.520 642.380 1402.500 729.380 ;
        RECT 315.520 552.380 1402.500 639.380 ;
        RECT 315.520 462.380 1402.500 549.380 ;
        RECT 315.520 395.670 1402.500 459.380 ;
      LAYER met5 ;
        RECT 315.520 319.080 1402.500 320.680 ;
        RECT 315.520 242.490 1402.500 244.090 ;
  END
END user_project_wrapper
END LIBRARY

