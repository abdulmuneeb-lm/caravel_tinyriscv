magic
tech sky130A
magscale 1 2
timestamp 1609742308
<< locali >>
rect 8125 685899 8159 695453
rect 72525 684607 72559 694093
rect 137845 685899 137879 695453
rect 219081 685899 219115 695453
rect 72801 676107 72835 684437
rect 154313 676243 154347 685797
rect 284033 676243 284067 685797
rect 218989 666587 219023 676141
rect 156613 40987 156647 41157
rect 270509 41123 270543 41293
rect 274741 41055 274775 41293
rect 280169 41055 280203 41157
rect 289737 41055 289771 41157
rect 331137 41157 331321 41191
rect 331137 41055 331171 41157
rect 289863 40953 289921 40987
rect 309149 40375 309183 40953
rect 338129 40919 338163 41157
rect 434821 29019 434855 38573
rect 383485 22015 383519 28917
rect 412649 19363 412683 26945
rect 372629 12291 372663 19261
rect 434821 9775 434855 19261
rect 395997 4675 396031 4777
rect 396089 4743 396123 4845
rect 405749 4743 405783 4845
rect 237297 3587 237331 3961
rect 132509 3315 132543 3485
rect 183385 3247 183419 3349
rect 365545 3043 365579 3553
rect 365637 3451 365671 3553
rect 412097 595 412131 9605
rect 413293 4675 413327 4845
rect 415685 595 415719 9605
rect 422953 4675 422987 4845
rect 427829 4675 427863 4845
rect 427771 4641 427863 4675
rect 435833 595 435867 9605
<< viali >>
rect 8125 695453 8159 695487
rect 137845 695453 137879 695487
rect 8125 685865 8159 685899
rect 72525 694093 72559 694127
rect 137845 685865 137879 685899
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 72525 684573 72559 684607
rect 154313 685797 154347 685831
rect 72801 684437 72835 684471
rect 154313 676209 154347 676243
rect 284033 685797 284067 685831
rect 284033 676209 284067 676243
rect 72801 676073 72835 676107
rect 218989 676141 219023 676175
rect 218989 666553 219023 666587
rect 270509 41293 270543 41327
rect 156613 41157 156647 41191
rect 270509 41089 270543 41123
rect 274741 41293 274775 41327
rect 274741 41021 274775 41055
rect 280169 41157 280203 41191
rect 280169 41021 280203 41055
rect 289737 41157 289771 41191
rect 289737 41021 289771 41055
rect 331321 41157 331355 41191
rect 338129 41157 338163 41191
rect 331137 41021 331171 41055
rect 156613 40953 156647 40987
rect 289829 40953 289863 40987
rect 289921 40953 289955 40987
rect 309149 40953 309183 40987
rect 338129 40885 338163 40919
rect 309149 40341 309183 40375
rect 434821 38573 434855 38607
rect 434821 28985 434855 29019
rect 383485 28917 383519 28951
rect 383485 21981 383519 22015
rect 412649 26945 412683 26979
rect 412649 19329 412683 19363
rect 372629 19261 372663 19295
rect 372629 12257 372663 12291
rect 434821 19261 434855 19295
rect 434821 9741 434855 9775
rect 412097 9605 412131 9639
rect 396089 4845 396123 4879
rect 395997 4777 396031 4811
rect 396089 4709 396123 4743
rect 405749 4845 405783 4879
rect 405749 4709 405783 4743
rect 395997 4641 396031 4675
rect 237297 3961 237331 3995
rect 237297 3553 237331 3587
rect 365545 3553 365579 3587
rect 132509 3485 132543 3519
rect 132509 3281 132543 3315
rect 183385 3349 183419 3383
rect 183385 3213 183419 3247
rect 365637 3553 365671 3587
rect 365637 3417 365671 3451
rect 365545 3009 365579 3043
rect 415685 9605 415719 9639
rect 413293 4845 413327 4879
rect 413293 4641 413327 4675
rect 412097 561 412131 595
rect 435833 9605 435867 9639
rect 422953 4845 422987 4879
rect 427829 4845 427863 4879
rect 422953 4641 422987 4675
rect 427737 4641 427771 4675
rect 415685 561 415719 595
rect 435833 561 435867 595
<< metal1 >>
rect 394602 700408 394608 700460
rect 394660 700448 394666 700460
rect 413646 700448 413652 700460
rect 394660 700420 413652 700448
rect 394660 700408 394666 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 463602 700408 463608 700460
rect 463660 700448 463666 700460
rect 494790 700448 494796 700460
rect 463660 700420 494796 700448
rect 463660 700408 463666 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 514662 700408 514668 700460
rect 514720 700448 514726 700460
rect 559650 700448 559656 700460
rect 514720 700420 559656 700448
rect 514720 700408 514726 700420
rect 559650 700408 559656 700420
rect 559708 700408 559714 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 411162 700340 411168 700392
rect 411220 700380 411226 700392
rect 429838 700380 429844 700392
rect 411220 700352 429844 700380
rect 411220 700340 411226 700352
rect 429838 700340 429844 700352
rect 429896 700340 429902 700392
rect 445662 700340 445668 700392
rect 445720 700380 445726 700392
rect 478506 700380 478512 700392
rect 445720 700352 478512 700380
rect 445720 700340 445726 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 496722 700340 496728 700392
rect 496780 700380 496786 700392
rect 543458 700380 543464 700392
rect 496780 700352 543464 700380
rect 496780 700340 496786 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 344278 700272 344284 700324
rect 344336 700312 344342 700324
rect 348786 700312 348792 700324
rect 344336 700284 348792 700312
rect 344336 700272 344342 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 378042 700272 378048 700324
rect 378100 700312 378106 700324
rect 397454 700312 397460 700324
rect 378100 700284 397460 700312
rect 378100 700272 378106 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 429102 700272 429108 700324
rect 429160 700312 429166 700324
rect 462314 700312 462320 700324
rect 429160 700284 462320 700312
rect 429160 700272 429166 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 480162 700272 480168 700324
rect 480220 700312 480226 700324
rect 527174 700312 527180 700324
rect 480220 700284 527180 700312
rect 480220 700272 480226 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 326982 699660 326988 699712
rect 327040 699700 327046 699712
rect 332502 699700 332508 699712
rect 327040 699672 332508 699700
rect 327040 699660 327046 699672
rect 332502 699660 332508 699672
rect 332560 699660 332566 699712
rect 360102 699660 360108 699712
rect 360160 699700 360166 699712
rect 364978 699700 364984 699712
rect 360160 699672 364984 699700
rect 360160 699660 360166 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 137738 698232 137744 698284
rect 137796 698272 137802 698284
rect 137922 698272 137928 698284
rect 137796 698244 137928 698272
rect 137796 698232 137802 698244
rect 137922 698232 137928 698244
rect 137980 698232 137986 698284
rect 523770 696940 523776 696992
rect 523828 696980 523834 696992
rect 580166 696980 580172 696992
rect 523828 696952 580172 696980
rect 523828 696940 523834 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 283834 695512 283840 695564
rect 283892 695552 283898 695564
rect 283926 695552 283932 695564
rect 283892 695524 283932 695552
rect 283892 695512 283898 695524
rect 283926 695512 283932 695524
rect 283984 695512 283990 695564
rect 8113 695487 8171 695493
rect 8113 695453 8125 695487
rect 8159 695484 8171 695487
rect 8202 695484 8208 695496
rect 8159 695456 8208 695484
rect 8159 695453 8171 695456
rect 8113 695447 8171 695453
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 137833 695487 137891 695493
rect 137833 695453 137845 695487
rect 137879 695484 137891 695487
rect 137922 695484 137928 695496
rect 137879 695456 137928 695484
rect 137879 695453 137891 695456
rect 137833 695447 137891 695453
rect 137922 695444 137928 695456
rect 137980 695444 137986 695496
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 72513 694127 72571 694133
rect 72513 694093 72525 694127
rect 72559 694124 72571 694127
rect 72694 694124 72700 694136
rect 72559 694096 72700 694124
rect 72559 694093 72571 694096
rect 72513 694087 72571 694093
rect 72694 694084 72700 694096
rect 72752 694084 72758 694136
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 283926 688576 283932 688628
rect 283984 688616 283990 688628
rect 284110 688616 284116 688628
rect 283984 688588 284116 688616
rect 283984 688576 283990 688588
rect 284110 688576 284116 688588
rect 284168 688576 284174 688628
rect 8110 685896 8116 685908
rect 8071 685868 8116 685896
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 137830 685896 137836 685908
rect 137791 685868 137836 685896
rect 137830 685856 137836 685868
rect 137888 685856 137894 685908
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 523678 685856 523684 685908
rect 523736 685896 523742 685908
rect 580166 685896 580172 685908
rect 523736 685868 580172 685896
rect 523736 685856 523742 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 284021 685831 284079 685837
rect 284021 685797 284033 685831
rect 284067 685828 284079 685831
rect 284110 685828 284116 685840
rect 284067 685800 284116 685828
rect 284067 685797 284079 685800
rect 284021 685791 284079 685797
rect 284110 685788 284116 685800
rect 284168 685788 284174 685840
rect 72510 684604 72516 684616
rect 72471 684576 72516 684604
rect 72510 684564 72516 684576
rect 72568 684564 72574 684616
rect 72510 684428 72516 684480
rect 72568 684468 72574 684480
rect 72789 684471 72847 684477
rect 72789 684468 72801 684471
rect 72568 684440 72801 684468
rect 72568 684428 72574 684440
rect 72789 684437 72801 684440
rect 72835 684437 72847 684471
rect 72789 684431 72847 684437
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 137830 679028 137836 679040
rect 137756 679000 137836 679028
rect 137756 678972 137784 679000
rect 137830 678988 137836 679000
rect 137888 678988 137894 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 137738 678920 137744 678972
rect 137796 678920 137802 678972
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 284018 676240 284024 676252
rect 283979 676212 284024 676240
rect 284018 676200 284024 676212
rect 284076 676200 284082 676252
rect 218974 676172 218980 676184
rect 218935 676144 218980 676172
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 72786 676104 72792 676116
rect 72747 676076 72792 676104
rect 72786 676064 72792 676076
rect 72844 676064 72850 676116
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 137738 673480 137744 673532
rect 137796 673520 137802 673532
rect 137922 673520 137928 673532
rect 137796 673492 137928 673520
rect 137796 673480 137802 673492
rect 137922 673480 137928 673492
rect 137980 673480 137986 673532
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 284018 673480 284024 673532
rect 284076 673520 284082 673532
rect 284202 673520 284208 673532
rect 284076 673492 284208 673520
rect 284076 673480 284082 673492
rect 284202 673480 284208 673492
rect 284260 673480 284266 673532
rect 72786 669332 72792 669384
rect 72844 669332 72850 669384
rect 72804 669248 72832 669332
rect 72786 669196 72792 669248
rect 72844 669196 72850 669248
rect 218977 666587 219035 666593
rect 218977 666553 218989 666587
rect 219023 666584 219035 666587
rect 219066 666584 219072 666596
rect 219023 666556 219072 666584
rect 219023 666553 219035 666556
rect 218977 666547 219035 666553
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 8018 654100 8024 654152
rect 8076 654140 8082 654152
rect 8202 654140 8208 654152
rect 8076 654112 8208 654140
rect 8076 654100 8082 654112
rect 8202 654100 8208 654112
rect 8260 654100 8266 654152
rect 137738 654100 137744 654152
rect 137796 654140 137802 654152
rect 137922 654140 137928 654152
rect 137796 654112 137928 654140
rect 137796 654100 137802 654112
rect 137922 654100 137928 654112
rect 137980 654100 137986 654152
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 284018 654100 284024 654152
rect 284076 654140 284082 654152
rect 284202 654140 284208 654152
rect 284076 654112 284208 654140
rect 284076 654100 284082 654112
rect 284202 654100 284208 654112
rect 284260 654100 284266 654152
rect 342990 645804 342996 645856
rect 343048 645844 343054 645856
rect 344278 645844 344284 645856
rect 343048 645816 344284 645844
rect 343048 645804 343054 645816
rect 344278 645804 344284 645816
rect 344336 645804 344342 645856
rect 377122 645804 377128 645856
rect 377180 645844 377186 645856
rect 378042 645844 378048 645856
rect 377180 645816 378048 645844
rect 377180 645804 377186 645816
rect 378042 645804 378048 645816
rect 378100 645804 378106 645856
rect 428182 645804 428188 645856
rect 428240 645844 428246 645856
rect 429102 645844 429108 645856
rect 428240 645816 429108 645844
rect 428240 645804 428246 645816
rect 429102 645804 429108 645816
rect 429160 645804 429166 645856
rect 462314 645804 462320 645856
rect 462372 645844 462378 645856
rect 463602 645844 463608 645856
rect 462372 645816 463608 645844
rect 462372 645804 462378 645816
rect 463602 645804 463608 645816
rect 463660 645804 463666 645856
rect 479334 645804 479340 645856
rect 479392 645844 479398 645856
rect 480162 645844 480168 645856
rect 479392 645816 480168 645844
rect 479392 645804 479398 645816
rect 480162 645804 480168 645816
rect 480220 645804 480226 645856
rect 513374 645600 513380 645652
rect 513432 645640 513438 645652
rect 514662 645640 514668 645652
rect 513432 645612 514668 645640
rect 513432 645600 513438 645612
rect 514662 645600 514668 645612
rect 514720 645600 514726 645652
rect 325970 645464 325976 645516
rect 326028 645504 326034 645516
rect 326982 645504 326988 645516
rect 326028 645476 326988 645504
rect 326028 645464 326034 645476
rect 326982 645464 326988 645476
rect 327040 645464 327046 645516
rect 73062 645328 73068 645380
rect 73120 645368 73126 645380
rect 121546 645368 121552 645380
rect 73120 645340 121552 645368
rect 73120 645328 73126 645340
rect 121546 645328 121552 645340
rect 121604 645328 121610 645380
rect 137922 645328 137928 645380
rect 137980 645368 137986 645380
rect 172698 645368 172704 645380
rect 137980 645340 172704 645368
rect 137980 645328 137986 645340
rect 172698 645328 172704 645340
rect 172756 645328 172762 645380
rect 8202 645260 8208 645312
rect 8260 645300 8266 645312
rect 70486 645300 70492 645312
rect 8260 645272 70492 645300
rect 8260 645260 8266 645272
rect 70486 645260 70492 645272
rect 70544 645260 70550 645312
rect 89622 645260 89628 645312
rect 89680 645300 89686 645312
rect 138566 645300 138572 645312
rect 89680 645272 138572 645300
rect 89680 645260 89686 645272
rect 138566 645260 138572 645272
rect 138624 645260 138630 645312
rect 41322 645192 41328 645244
rect 41380 645232 41386 645244
rect 104526 645232 104532 645244
rect 41380 645204 104532 645232
rect 41380 645192 41386 645204
rect 104526 645192 104532 645204
rect 104584 645192 104590 645244
rect 154482 645192 154488 645244
rect 154540 645232 154546 645244
rect 189718 645232 189724 645244
rect 154540 645204 189724 645232
rect 154540 645192 154546 645204
rect 189718 645192 189724 645204
rect 189776 645192 189782 645244
rect 202782 645192 202788 645244
rect 202840 645232 202846 645244
rect 223758 645232 223764 645244
rect 202840 645204 223764 645232
rect 202840 645192 202846 645204
rect 223758 645192 223764 645204
rect 223816 645192 223822 645244
rect 235902 645192 235908 645244
rect 235960 645232 235966 645244
rect 257890 645232 257896 645244
rect 235960 645204 257896 645232
rect 235960 645192 235966 645204
rect 257890 645192 257896 645204
rect 257948 645192 257954 645244
rect 24762 645124 24768 645176
rect 24820 645164 24826 645176
rect 87506 645164 87512 645176
rect 24820 645136 87512 645164
rect 24820 645124 24826 645136
rect 87506 645124 87512 645136
rect 87564 645124 87570 645176
rect 106182 645124 106188 645176
rect 106240 645164 106246 645176
rect 155586 645164 155592 645176
rect 106240 645136 155592 645164
rect 106240 645124 106246 645136
rect 155586 645124 155592 645136
rect 155644 645124 155650 645176
rect 171042 645124 171048 645176
rect 171100 645164 171106 645176
rect 206738 645164 206744 645176
rect 171100 645136 206744 645164
rect 171100 645124 171106 645136
rect 206738 645124 206744 645136
rect 206796 645124 206802 645176
rect 219342 645124 219348 645176
rect 219400 645164 219406 645176
rect 240778 645164 240784 645176
rect 219400 645136 240784 645164
rect 219400 645124 219406 645136
rect 240778 645124 240784 645136
rect 240836 645124 240842 645176
rect 267642 645124 267648 645176
rect 267700 645164 267706 645176
rect 274910 645164 274916 645176
rect 267700 645136 274916 645164
rect 267700 645124 267706 645136
rect 274910 645124 274916 645136
rect 274968 645124 274974 645176
rect 284202 645124 284208 645176
rect 284260 645164 284266 645176
rect 291930 645164 291936 645176
rect 284260 645136 291936 645164
rect 284260 645124 284266 645136
rect 291930 645124 291936 645136
rect 291988 645124 291994 645176
rect 300762 644852 300768 644904
rect 300820 644892 300826 644904
rect 308950 644892 308956 644904
rect 300820 644864 308956 644892
rect 300820 644852 300826 644864
rect 308950 644852 308956 644864
rect 309008 644852 309014 644904
rect 523862 638936 523868 638988
rect 523920 638976 523926 638988
rect 580166 638976 580172 638988
rect 523920 638948 580172 638976
rect 523920 638936 523926 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 3418 636148 3424 636200
rect 3476 636188 3482 636200
rect 59354 636188 59360 636200
rect 3476 636160 59360 636188
rect 3476 636148 3482 636160
rect 59354 636148 59360 636160
rect 59412 636148 59418 636200
rect 3510 622344 3516 622396
rect 3568 622384 3574 622396
rect 59354 622384 59360 622396
rect 3568 622356 59360 622384
rect 3568 622344 3574 622356
rect 59354 622344 59360 622356
rect 59412 622344 59418 622396
rect 524322 609900 524328 609952
rect 524380 609940 524386 609952
rect 580258 609940 580264 609952
rect 524380 609912 580264 609940
rect 524380 609900 524386 609912
rect 580258 609900 580264 609912
rect 580316 609900 580322 609952
rect 3602 608540 3608 608592
rect 3660 608580 3666 608592
rect 59354 608580 59360 608592
rect 3660 608552 59360 608580
rect 3660 608540 3666 608552
rect 59354 608540 59360 608552
rect 59412 608540 59418 608592
rect 523770 603100 523776 603152
rect 523828 603140 523834 603152
rect 580166 603140 580172 603152
rect 523828 603112 580172 603140
rect 523828 603100 523834 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 523678 597456 523684 597508
rect 523736 597496 523742 597508
rect 580442 597496 580448 597508
rect 523736 597468 580448 597496
rect 523736 597456 523742 597468
rect 580442 597456 580448 597468
rect 580500 597456 580506 597508
rect 3418 593308 3424 593360
rect 3476 593348 3482 593360
rect 59354 593348 59360 593360
rect 3476 593320 59360 593348
rect 3476 593308 3482 593320
rect 59354 593308 59360 593320
rect 59412 593308 59418 593360
rect 523678 592016 523684 592068
rect 523736 592056 523742 592068
rect 580166 592056 580172 592068
rect 523736 592028 580172 592056
rect 523736 592016 523742 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 3510 579572 3516 579624
rect 3568 579612 3574 579624
rect 59354 579612 59360 579624
rect 3568 579584 59360 579612
rect 3568 579572 3574 579584
rect 59354 579572 59360 579584
rect 59412 579572 59418 579624
rect 524322 569848 524328 569900
rect 524380 569888 524386 569900
rect 580350 569888 580356 569900
rect 524380 569860 580356 569888
rect 524380 569848 524386 569860
rect 580350 569848 580356 569860
rect 580408 569848 580414 569900
rect 3602 565768 3608 565820
rect 3660 565808 3666 565820
rect 59354 565808 59360 565820
rect 3660 565780 59360 565808
rect 3660 565768 3666 565780
rect 59354 565768 59360 565780
rect 59412 565768 59418 565820
rect 523862 556180 523868 556232
rect 523920 556220 523926 556232
rect 580166 556220 580172 556232
rect 523920 556192 580172 556220
rect 523920 556180 523926 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 3418 550536 3424 550588
rect 3476 550576 3482 550588
rect 59354 550576 59360 550588
rect 3476 550548 59360 550576
rect 3476 550536 3482 550548
rect 59354 550536 59360 550548
rect 59412 550536 59418 550588
rect 523770 545096 523776 545148
rect 523828 545136 523834 545148
rect 580166 545136 580172 545148
rect 523828 545108 580172 545136
rect 523828 545096 523834 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 3510 536732 3516 536784
rect 3568 536772 3574 536784
rect 59354 536772 59360 536784
rect 3568 536744 59360 536772
rect 3568 536732 3574 536744
rect 59354 536732 59360 536744
rect 59412 536732 59418 536784
rect 523218 531224 523224 531276
rect 523276 531264 523282 531276
rect 580258 531264 580264 531276
rect 523276 531236 580264 531264
rect 523276 531224 523282 531236
rect 580258 531224 580264 531236
rect 580316 531224 580322 531276
rect 3418 522928 3424 522980
rect 3476 522968 3482 522980
rect 59354 522968 59360 522980
rect 3476 522940 59360 522968
rect 3476 522928 3482 522940
rect 59354 522928 59360 522940
rect 59412 522928 59418 522980
rect 523862 509260 523868 509312
rect 523920 509300 523926 509312
rect 580166 509300 580172 509312
rect 523920 509272 580172 509300
rect 523920 509260 523926 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 3326 507764 3332 507816
rect 3384 507804 3390 507816
rect 59354 507804 59360 507816
rect 3384 507776 59360 507804
rect 3384 507764 3390 507776
rect 59354 507764 59360 507776
rect 59412 507764 59418 507816
rect 523770 498176 523776 498228
rect 523828 498216 523834 498228
rect 580166 498216 580172 498228
rect 523828 498188 580172 498216
rect 523828 498176 523834 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 3326 493960 3332 494012
rect 3384 494000 3390 494012
rect 59354 494000 59360 494012
rect 3384 493972 59360 494000
rect 3384 493960 3390 493972
rect 59354 493960 59360 493972
rect 59412 493960 59418 494012
rect 524322 491240 524328 491292
rect 524380 491280 524386 491292
rect 580350 491280 580356 491292
rect 524380 491252 580356 491280
rect 524380 491240 524386 491252
rect 580350 491240 580356 491252
rect 580408 491240 580414 491292
rect 523678 485800 523684 485852
rect 523736 485840 523742 485852
rect 580166 485840 580172 485852
rect 523736 485812 580172 485840
rect 523736 485800 523742 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 3602 480156 3608 480208
rect 3660 480196 3666 480208
rect 59354 480196 59360 480208
rect 3660 480168 59360 480196
rect 3660 480156 3666 480168
rect 59354 480156 59360 480168
rect 59412 480156 59418 480208
rect 3418 463700 3424 463752
rect 3476 463740 3482 463752
rect 59354 463740 59360 463752
rect 3476 463712 59360 463740
rect 3476 463700 3482 463712
rect 59354 463700 59360 463712
rect 59412 463700 59418 463752
rect 523862 462340 523868 462392
rect 523920 462380 523926 462392
rect 580166 462380 580172 462392
rect 523920 462352 580172 462380
rect 523920 462340 523926 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 523770 451256 523776 451308
rect 523828 451296 523834 451308
rect 580166 451296 580172 451308
rect 523828 451268 580172 451296
rect 523828 451256 523834 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 3418 449896 3424 449948
rect 3476 449936 3482 449948
rect 59354 449936 59360 449948
rect 3476 449908 59360 449936
rect 3476 449896 3482 449908
rect 59354 449896 59360 449908
rect 59412 449896 59418 449948
rect 523678 438880 523684 438932
rect 523736 438920 523742 438932
rect 580166 438920 580172 438932
rect 523736 438892 580172 438920
rect 523736 438880 523742 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 3418 436092 3424 436144
rect 3476 436132 3482 436144
rect 59354 436132 59360 436144
rect 3476 436104 59360 436132
rect 3476 436092 3482 436104
rect 59354 436092 59360 436104
rect 59412 436092 59418 436144
rect 3510 420928 3516 420980
rect 3568 420968 3574 420980
rect 59354 420968 59360 420980
rect 3568 420940 59360 420968
rect 3568 420928 3574 420940
rect 59354 420928 59360 420940
rect 59412 420928 59418 420980
rect 523862 415420 523868 415472
rect 523920 415460 523926 415472
rect 580166 415460 580172 415472
rect 523920 415432 580172 415460
rect 523920 415420 523926 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 3418 407124 3424 407176
rect 3476 407164 3482 407176
rect 59354 407164 59360 407176
rect 3476 407136 59360 407164
rect 3476 407124 3482 407136
rect 59354 407124 59360 407136
rect 59412 407124 59418 407176
rect 523770 404336 523776 404388
rect 523828 404376 523834 404388
rect 580166 404376 580172 404388
rect 523828 404348 580172 404376
rect 523828 404336 523834 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 391960 3516 392012
rect 3568 392000 3574 392012
rect 59354 392000 59360 392012
rect 3568 391972 59360 392000
rect 3568 391960 3574 391972
rect 59354 391960 59360 391972
rect 59412 391960 59418 392012
rect 523678 391960 523684 392012
rect 523736 392000 523742 392012
rect 580166 392000 580172 392012
rect 523736 391972 580172 392000
rect 523736 391960 523742 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 3418 378156 3424 378208
rect 3476 378196 3482 378208
rect 59354 378196 59360 378208
rect 3476 378168 59360 378196
rect 3476 378156 3482 378168
rect 59354 378156 59360 378168
rect 59412 378156 59418 378208
rect 523678 368500 523684 368552
rect 523736 368540 523742 368552
rect 580166 368540 580172 368552
rect 523736 368512 580172 368540
rect 523736 368500 523742 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 3510 364352 3516 364404
rect 3568 364392 3574 364404
rect 59354 364392 59360 364404
rect 3568 364364 59360 364392
rect 3568 364352 3574 364364
rect 59354 364352 59360 364364
rect 59412 364352 59418 364404
rect 523770 357416 523776 357468
rect 523828 357456 523834 357468
rect 580166 357456 580172 357468
rect 523828 357428 580172 357456
rect 523828 357416 523834 357428
rect 580166 357416 580172 357428
rect 580224 357416 580230 357468
rect 3602 349120 3608 349172
rect 3660 349160 3666 349172
rect 59354 349160 59360 349172
rect 3660 349132 59360 349160
rect 3660 349120 3666 349132
rect 59354 349120 59360 349132
rect 59412 349120 59418 349172
rect 523678 345040 523684 345092
rect 523736 345080 523742 345092
rect 580166 345080 580172 345092
rect 523736 345052 580172 345080
rect 523736 345040 523742 345052
rect 580166 345040 580172 345052
rect 580224 345040 580230 345092
rect 3418 335316 3424 335368
rect 3476 335356 3482 335368
rect 59354 335356 59360 335368
rect 3476 335328 59360 335356
rect 3476 335316 3482 335328
rect 59354 335316 59360 335328
rect 59412 335316 59418 335368
rect 3510 321580 3516 321632
rect 3568 321620 3574 321632
rect 59354 321620 59360 321632
rect 3568 321592 59360 321620
rect 3568 321580 3574 321592
rect 59354 321580 59360 321592
rect 59412 321580 59418 321632
rect 523494 321580 523500 321632
rect 523552 321620 523558 321632
rect 580166 321620 580172 321632
rect 523552 321592 580172 321620
rect 523552 321580 523558 321592
rect 580166 321580 580172 321592
rect 580224 321580 580230 321632
rect 523678 310496 523684 310548
rect 523736 310536 523742 310548
rect 579798 310536 579804 310548
rect 523736 310508 579804 310536
rect 523736 310496 523742 310508
rect 579798 310496 579804 310508
rect 579856 310496 579862 310548
rect 3694 306348 3700 306400
rect 3752 306388 3758 306400
rect 59354 306388 59360 306400
rect 3752 306360 59360 306388
rect 3752 306348 3758 306360
rect 59354 306348 59360 306360
rect 59412 306348 59418 306400
rect 523218 298120 523224 298172
rect 523276 298160 523282 298172
rect 580166 298160 580172 298172
rect 523276 298132 580172 298160
rect 523276 298120 523282 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3602 292544 3608 292596
rect 3660 292584 3666 292596
rect 59354 292584 59360 292596
rect 3660 292556 59360 292584
rect 3660 292544 3666 292556
rect 59354 292544 59360 292556
rect 59412 292544 59418 292596
rect 3418 278740 3424 278792
rect 3476 278780 3482 278792
rect 59354 278780 59360 278792
rect 3476 278752 59360 278780
rect 3476 278740 3482 278752
rect 59354 278740 59360 278752
rect 59412 278740 59418 278792
rect 524322 275952 524328 276004
rect 524380 275992 524386 276004
rect 580166 275992 580172 276004
rect 524380 275964 580172 275992
rect 524380 275952 524386 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 3694 263576 3700 263628
rect 3752 263616 3758 263628
rect 59354 263616 59360 263628
rect 3752 263588 59360 263616
rect 3752 263576 3758 263588
rect 59354 263576 59360 263588
rect 59412 263576 59418 263628
rect 524322 263576 524328 263628
rect 524380 263616 524386 263628
rect 579798 263616 579804 263628
rect 524380 263588 579804 263616
rect 524380 263576 524386 263588
rect 579798 263576 579804 263588
rect 579856 263576 579862 263628
rect 523954 251200 523960 251252
rect 524012 251240 524018 251252
rect 580166 251240 580172 251252
rect 524012 251212 580172 251240
rect 524012 251200 524018 251212
rect 580166 251200 580172 251212
rect 580224 251200 580230 251252
rect 3510 249772 3516 249824
rect 3568 249812 3574 249824
rect 59354 249812 59360 249824
rect 3568 249784 59360 249812
rect 3568 249772 3574 249784
rect 59354 249772 59360 249784
rect 59412 249772 59418 249824
rect 3602 235968 3608 236020
rect 3660 236008 3666 236020
rect 59354 236008 59360 236020
rect 3660 235980 59360 236008
rect 3660 235968 3666 235980
rect 59354 235968 59360 235980
rect 59412 235968 59418 236020
rect 523678 229032 523684 229084
rect 523736 229072 523742 229084
rect 580166 229072 580172 229084
rect 523736 229044 580172 229072
rect 523736 229032 523742 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 3418 220804 3424 220856
rect 3476 220844 3482 220856
rect 59354 220844 59360 220856
rect 3476 220816 59360 220844
rect 3476 220804 3482 220816
rect 59354 220804 59360 220816
rect 59412 220804 59418 220856
rect 523678 217948 523684 218000
rect 523736 217988 523742 218000
rect 580166 217988 580172 218000
rect 523736 217960 580172 217988
rect 523736 217948 523742 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 3694 207000 3700 207052
rect 3752 207040 3758 207052
rect 59354 207040 59360 207052
rect 3752 207012 59360 207040
rect 3752 207000 3758 207012
rect 59354 207000 59360 207012
rect 59412 207000 59418 207052
rect 523402 205572 523408 205624
rect 523460 205612 523466 205624
rect 579798 205612 579804 205624
rect 523460 205584 579804 205612
rect 523460 205572 523466 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 3602 191836 3608 191888
rect 3660 191876 3666 191888
rect 59354 191876 59360 191888
rect 3660 191848 59360 191876
rect 3660 191836 3666 191848
rect 59354 191836 59360 191848
rect 59412 191836 59418 191888
rect 523678 182112 523684 182164
rect 523736 182152 523742 182164
rect 580166 182152 580172 182164
rect 523736 182124 580172 182152
rect 523736 182112 523742 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 3510 178032 3516 178084
rect 3568 178072 3574 178084
rect 59354 178072 59360 178084
rect 3568 178044 59360 178072
rect 3568 178032 3574 178044
rect 59354 178032 59360 178044
rect 59412 178032 59418 178084
rect 523770 171028 523776 171080
rect 523828 171068 523834 171080
rect 580166 171068 580172 171080
rect 523828 171040 580172 171068
rect 523828 171028 523834 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 3418 164228 3424 164280
rect 3476 164268 3482 164280
rect 59354 164268 59360 164280
rect 3476 164240 59360 164268
rect 3476 164228 3482 164240
rect 59354 164228 59360 164240
rect 59412 164228 59418 164280
rect 523678 158652 523684 158704
rect 523736 158692 523742 158704
rect 579798 158692 579804 158704
rect 523736 158664 579804 158692
rect 523736 158652 523742 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 3694 149064 3700 149116
rect 3752 149104 3758 149116
rect 59354 149104 59360 149116
rect 3752 149076 59360 149104
rect 3752 149064 3758 149076
rect 59354 149064 59360 149076
rect 59412 149064 59418 149116
rect 3602 135260 3608 135312
rect 3660 135300 3666 135312
rect 59354 135300 59360 135312
rect 3660 135272 59360 135300
rect 3660 135260 3666 135272
rect 59354 135260 59360 135272
rect 59412 135260 59418 135312
rect 523678 135192 523684 135244
rect 523736 135232 523742 135244
rect 580166 135232 580172 135244
rect 523736 135204 580172 135232
rect 523736 135192 523742 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 523862 124108 523868 124160
rect 523920 124148 523926 124160
rect 580166 124148 580172 124160
rect 523920 124120 580172 124148
rect 523920 124108 523926 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 3510 121456 3516 121508
rect 3568 121496 3574 121508
rect 59354 121496 59360 121508
rect 3568 121468 59360 121496
rect 3568 121456 3574 121468
rect 59354 121456 59360 121468
rect 59412 121456 59418 121508
rect 523770 111732 523776 111784
rect 523828 111772 523834 111784
rect 579798 111772 579804 111784
rect 523828 111744 579804 111772
rect 523828 111732 523834 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 3786 106292 3792 106344
rect 3844 106332 3850 106344
rect 59354 106332 59360 106344
rect 3844 106304 59360 106332
rect 3844 106292 3850 106304
rect 59354 106292 59360 106304
rect 59412 106292 59418 106344
rect 3694 92488 3700 92540
rect 3752 92528 3758 92540
rect 59354 92528 59360 92540
rect 3752 92500 59360 92528
rect 3752 92488 3758 92500
rect 59354 92488 59360 92500
rect 59412 92488 59418 92540
rect 523678 88272 523684 88324
rect 523736 88312 523742 88324
rect 580166 88312 580172 88324
rect 523736 88284 580172 88312
rect 523736 88272 523742 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 3418 78684 3424 78736
rect 3476 78724 3482 78736
rect 59354 78724 59360 78736
rect 3476 78696 59360 78724
rect 3476 78684 3482 78696
rect 59354 78684 59360 78696
rect 59412 78684 59418 78736
rect 523770 77188 523776 77240
rect 523828 77228 523834 77240
rect 580166 77228 580172 77240
rect 523828 77200 580172 77228
rect 523828 77188 523834 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 523862 64812 523868 64864
rect 523920 64852 523926 64864
rect 579798 64852 579804 64864
rect 523920 64824 579804 64852
rect 523920 64812 523926 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 3602 63520 3608 63572
rect 3660 63560 3666 63572
rect 59354 63560 59360 63572
rect 3660 63532 59360 63560
rect 3660 63520 3666 63532
rect 59354 63520 59360 63532
rect 59412 63520 59418 63572
rect 3510 49716 3516 49768
rect 3568 49756 3574 49768
rect 59354 49756 59360 49768
rect 3568 49728 59360 49756
rect 3568 49716 3574 49728
rect 59354 49716 59360 49728
rect 59412 49716 59418 49768
rect 523678 41352 523684 41404
rect 523736 41392 523742 41404
rect 580166 41392 580172 41404
rect 523736 41364 580172 41392
rect 523736 41352 523742 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 270497 41327 270555 41333
rect 270497 41293 270509 41327
rect 270543 41324 270555 41327
rect 274729 41327 274787 41333
rect 274729 41324 274741 41327
rect 270543 41296 274741 41324
rect 270543 41293 270555 41296
rect 270497 41287 270555 41293
rect 274729 41293 274741 41296
rect 274775 41293 274787 41327
rect 274729 41287 274787 41293
rect 272242 41216 272248 41268
rect 272300 41256 272306 41268
rect 273162 41256 273168 41268
rect 272300 41228 273168 41256
rect 272300 41216 272306 41228
rect 273162 41216 273168 41228
rect 273220 41216 273226 41268
rect 369946 41216 369952 41268
rect 370004 41256 370010 41268
rect 371050 41256 371056 41268
rect 370004 41228 371056 41256
rect 370004 41216 370010 41228
rect 371050 41216 371056 41228
rect 371108 41216 371114 41268
rect 145926 41148 145932 41200
rect 145984 41188 145990 41200
rect 156601 41191 156659 41197
rect 156601 41188 156613 41191
rect 145984 41160 156613 41188
rect 145984 41148 145990 41160
rect 156601 41157 156613 41160
rect 156647 41157 156659 41191
rect 156601 41151 156659 41157
rect 167362 41148 167368 41200
rect 167420 41188 167426 41200
rect 227898 41188 227904 41200
rect 167420 41160 227904 41188
rect 167420 41148 167426 41160
rect 227898 41148 227904 41160
rect 227956 41148 227962 41200
rect 253198 41148 253204 41200
rect 253256 41188 253262 41200
rect 280157 41191 280215 41197
rect 253256 41160 253980 41188
rect 253256 41148 253262 41160
rect 110230 41080 110236 41132
rect 110288 41120 110294 41132
rect 171226 41120 171232 41132
rect 110288 41092 171232 41120
rect 110288 41080 110294 41092
rect 171226 41080 171232 41092
rect 171284 41080 171290 41132
rect 188890 41080 188896 41132
rect 188948 41120 188954 41132
rect 249886 41120 249892 41132
rect 188948 41092 249892 41120
rect 188948 41080 188954 41092
rect 249886 41080 249892 41092
rect 249944 41080 249950 41132
rect 253952 41120 253980 41160
rect 280157 41157 280169 41191
rect 280203 41188 280215 41191
rect 289725 41191 289783 41197
rect 289725 41188 289737 41191
rect 280203 41160 289737 41188
rect 280203 41157 280215 41160
rect 280157 41151 280215 41157
rect 289725 41157 289737 41160
rect 289771 41157 289783 41191
rect 289725 41151 289783 41157
rect 331309 41191 331367 41197
rect 331309 41157 331321 41191
rect 331355 41188 331367 41191
rect 338117 41191 338175 41197
rect 338117 41188 338129 41191
rect 331355 41160 338129 41188
rect 331355 41157 331367 41160
rect 331309 41151 331367 41157
rect 338117 41157 338129 41160
rect 338163 41157 338175 41191
rect 338117 41151 338175 41157
rect 270497 41123 270555 41129
rect 270497 41120 270509 41123
rect 253952 41092 270509 41120
rect 270497 41089 270509 41092
rect 270543 41089 270555 41123
rect 270497 41083 270555 41089
rect 396166 41080 396172 41132
rect 396224 41120 396230 41132
rect 456886 41120 456892 41132
rect 396224 41092 456892 41120
rect 396224 41080 396230 41092
rect 456886 41080 456892 41092
rect 456944 41080 456950 41132
rect 131666 41012 131672 41064
rect 131724 41052 131730 41064
rect 193398 41052 193404 41064
rect 131724 41024 193404 41052
rect 131724 41012 131730 41024
rect 193398 41012 193404 41024
rect 193456 41012 193462 41064
rect 274729 41055 274787 41061
rect 274729 41021 274741 41055
rect 274775 41052 274787 41055
rect 280157 41055 280215 41061
rect 280157 41052 280169 41055
rect 274775 41024 280169 41052
rect 274775 41021 274787 41024
rect 274729 41015 274787 41021
rect 280157 41021 280169 41024
rect 280203 41021 280215 41055
rect 280157 41015 280215 41021
rect 289725 41055 289783 41061
rect 289725 41021 289737 41055
rect 289771 41052 289783 41055
rect 289771 41024 289860 41052
rect 289771 41021 289783 41024
rect 289725 41015 289783 41021
rect 81618 40944 81624 40996
rect 81676 40984 81682 40996
rect 142246 40984 142252 40996
rect 81676 40956 142252 40984
rect 81676 40944 81682 40956
rect 142246 40944 142252 40956
rect 142304 40944 142310 40996
rect 156601 40987 156659 40993
rect 156601 40953 156613 40987
rect 156647 40984 156659 40987
rect 207106 40984 207112 40996
rect 156647 40956 207112 40984
rect 156647 40953 156659 40956
rect 156601 40947 156659 40953
rect 207106 40944 207112 40956
rect 207164 40944 207170 40996
rect 210326 40944 210332 40996
rect 210384 40984 210390 40996
rect 270494 40984 270500 40996
rect 210384 40956 270500 40984
rect 210384 40944 210390 40956
rect 270494 40944 270500 40956
rect 270552 40944 270558 40996
rect 289832 40993 289860 41024
rect 318702 41012 318708 41064
rect 318760 41052 318766 41064
rect 331125 41055 331183 41061
rect 331125 41052 331137 41055
rect 318760 41024 331137 41052
rect 318760 41012 318766 41024
rect 331125 41021 331137 41024
rect 331171 41021 331183 41055
rect 331125 41015 331183 41021
rect 343726 41012 343732 41064
rect 343784 41052 343790 41064
rect 344830 41052 344836 41064
rect 343784 41024 344836 41052
rect 343784 41012 343790 41024
rect 344830 41012 344836 41024
rect 344888 41012 344894 41064
rect 367646 41012 367652 41064
rect 367704 41052 367710 41064
rect 367704 41024 369900 41052
rect 367704 41012 367710 41024
rect 289817 40987 289875 40993
rect 289817 40953 289829 40987
rect 289863 40953 289875 40987
rect 289817 40947 289875 40953
rect 289909 40987 289967 40993
rect 289909 40953 289921 40987
rect 289955 40984 289967 40987
rect 309137 40987 309195 40993
rect 309137 40984 309149 40987
rect 289955 40956 309149 40984
rect 289955 40953 289967 40956
rect 289909 40947 289967 40953
rect 309137 40953 309149 40956
rect 309183 40953 309195 40987
rect 369872 40984 369900 41024
rect 403342 41012 403348 41064
rect 403400 41052 403406 41064
rect 463786 41052 463792 41064
rect 403400 41024 463792 41052
rect 403400 41012 403406 41024
rect 463786 41012 463792 41024
rect 463844 41012 463850 41064
rect 427906 40984 427912 40996
rect 369872 40956 427912 40984
rect 309137 40947 309195 40953
rect 427906 40944 427912 40956
rect 427964 40944 427970 40996
rect 103054 40876 103060 40928
rect 103112 40916 103118 40928
rect 164326 40916 164332 40928
rect 103112 40888 164332 40916
rect 103112 40876 103118 40888
rect 164326 40876 164332 40888
rect 164384 40876 164390 40928
rect 174538 40876 174544 40928
rect 174596 40916 174602 40928
rect 236178 40916 236184 40928
rect 174596 40888 236184 40916
rect 174596 40876 174602 40888
rect 236178 40876 236184 40888
rect 236236 40876 236242 40928
rect 267642 40876 267648 40928
rect 267700 40916 267706 40928
rect 328546 40916 328552 40928
rect 267700 40888 328552 40916
rect 267700 40876 267706 40888
rect 328546 40876 328552 40888
rect 328604 40876 328610 40928
rect 338117 40919 338175 40925
rect 338117 40885 338129 40919
rect 338163 40916 338175 40919
rect 345658 40916 345664 40928
rect 338163 40888 345664 40916
rect 338163 40885 338175 40888
rect 338117 40879 338175 40885
rect 345658 40876 345664 40888
rect 345716 40876 345722 40928
rect 374730 40876 374736 40928
rect 374788 40916 374794 40928
rect 434806 40916 434812 40928
rect 374788 40888 434812 40916
rect 374788 40876 374794 40888
rect 434806 40876 434812 40888
rect 434864 40876 434870 40928
rect 474826 40876 474832 40928
rect 474884 40916 474890 40928
rect 535454 40916 535460 40928
rect 474884 40888 535460 40916
rect 474884 40876 474890 40888
rect 535454 40876 535460 40888
rect 535512 40876 535518 40928
rect 95878 40808 95884 40860
rect 95936 40848 95942 40860
rect 157426 40848 157432 40860
rect 95936 40820 157432 40848
rect 95936 40808 95942 40820
rect 157426 40808 157432 40820
rect 157484 40808 157490 40860
rect 181714 40808 181720 40860
rect 181772 40848 181778 40860
rect 242986 40848 242992 40860
rect 181772 40820 242992 40848
rect 181772 40808 181778 40820
rect 242986 40808 242992 40820
rect 243044 40808 243050 40860
rect 260374 40808 260380 40860
rect 260432 40848 260438 40860
rect 321738 40848 321744 40860
rect 260432 40820 321744 40848
rect 260432 40808 260438 40820
rect 321738 40808 321744 40820
rect 321796 40808 321802 40860
rect 381906 40808 381912 40860
rect 381964 40848 381970 40860
rect 443178 40848 443184 40860
rect 381964 40820 443184 40848
rect 381964 40808 381970 40820
rect 443178 40808 443184 40820
rect 443236 40808 443242 40860
rect 489178 40808 489184 40860
rect 489236 40848 489242 40860
rect 549254 40848 549260 40860
rect 489236 40820 549260 40848
rect 489236 40808 489242 40820
rect 549254 40808 549260 40820
rect 549312 40808 549318 40860
rect 88702 40740 88708 40792
rect 88760 40780 88766 40792
rect 150618 40780 150624 40792
rect 88760 40752 150624 40780
rect 88760 40740 88766 40752
rect 150618 40740 150624 40752
rect 150676 40740 150682 40792
rect 224586 40740 224592 40792
rect 224644 40780 224650 40792
rect 285766 40780 285772 40792
rect 224644 40752 285772 40780
rect 224644 40740 224650 40752
rect 285766 40740 285772 40752
rect 285824 40740 285830 40792
rect 333054 40740 333060 40792
rect 333112 40780 333118 40792
rect 333882 40780 333888 40792
rect 333112 40752 333888 40780
rect 333112 40740 333118 40752
rect 333882 40740 333888 40752
rect 333940 40740 333946 40792
rect 334250 40740 334256 40792
rect 334308 40780 334314 40792
rect 367738 40780 367744 40792
rect 334308 40752 367744 40780
rect 334308 40740 334314 40752
rect 367738 40740 367744 40752
rect 367796 40740 367802 40792
rect 389082 40740 389088 40792
rect 389140 40780 389146 40792
rect 449986 40780 449992 40792
rect 389140 40752 449992 40780
rect 389140 40740 389146 40752
rect 449986 40740 449992 40752
rect 450044 40740 450050 40792
rect 459370 40740 459376 40792
rect 459428 40780 459434 40792
rect 467098 40780 467104 40792
rect 459428 40752 467104 40780
rect 459428 40740 459434 40752
rect 467098 40740 467104 40752
rect 467156 40740 467162 40792
rect 482002 40740 482008 40792
rect 482060 40780 482066 40792
rect 542354 40780 542360 40792
rect 482060 40752 542360 40780
rect 482060 40740 482066 40752
rect 542354 40740 542360 40752
rect 542412 40740 542418 40792
rect 2682 40672 2688 40724
rect 2740 40712 2746 40724
rect 63678 40712 63684 40724
rect 2740 40684 63684 40712
rect 2740 40672 2746 40684
rect 63678 40672 63684 40684
rect 63736 40672 63742 40724
rect 67266 40672 67272 40724
rect 67324 40712 67330 40724
rect 128446 40712 128452 40724
rect 67324 40684 128452 40712
rect 67324 40672 67330 40684
rect 128446 40672 128452 40684
rect 128504 40672 128510 40724
rect 138842 40672 138848 40724
rect 138900 40712 138906 40724
rect 200206 40712 200212 40724
rect 138900 40684 200212 40712
rect 138900 40672 138906 40684
rect 200206 40672 200212 40684
rect 200264 40672 200270 40724
rect 217410 40672 217416 40724
rect 217468 40712 217474 40724
rect 278958 40712 278964 40724
rect 217468 40684 278964 40712
rect 217468 40672 217474 40684
rect 278958 40672 278964 40684
rect 279016 40672 279022 40724
rect 316402 40672 316408 40724
rect 316460 40712 316466 40724
rect 317322 40712 317328 40724
rect 316460 40684 317328 40712
rect 316460 40672 316466 40684
rect 317322 40672 317328 40684
rect 317380 40672 317386 40724
rect 324682 40672 324688 40724
rect 324740 40712 324746 40724
rect 325602 40712 325608 40724
rect 324740 40684 325608 40712
rect 324740 40672 324746 40684
rect 325602 40672 325608 40684
rect 325660 40672 325666 40724
rect 346118 40672 346124 40724
rect 346176 40712 346182 40724
rect 407206 40712 407212 40724
rect 346176 40684 407212 40712
rect 346176 40672 346182 40684
rect 407206 40672 407212 40684
rect 407264 40672 407270 40724
rect 467742 40672 467748 40724
rect 467800 40712 467806 40724
rect 528554 40712 528560 40724
rect 467800 40684 528560 40712
rect 467800 40672 467806 40684
rect 528554 40672 528560 40684
rect 528612 40672 528618 40724
rect 378318 40604 378324 40656
rect 378376 40644 378382 40656
rect 379422 40644 379428 40656
rect 378376 40616 379428 40644
rect 378376 40604 378382 40616
rect 379422 40604 379428 40616
rect 379480 40604 379486 40656
rect 247218 40536 247224 40588
rect 247276 40576 247282 40588
rect 248322 40576 248328 40588
rect 247276 40548 248328 40576
rect 247276 40536 247282 40548
rect 248322 40536 248328 40548
rect 248380 40536 248386 40588
rect 299658 40536 299664 40588
rect 299716 40576 299722 40588
rect 300762 40576 300768 40588
rect 299716 40548 300768 40576
rect 299716 40536 299722 40548
rect 300762 40536 300768 40548
rect 300820 40536 300826 40588
rect 290182 40468 290188 40520
rect 290240 40508 290246 40520
rect 291102 40508 291108 40520
rect 290240 40480 291108 40508
rect 290240 40468 290246 40480
rect 291102 40468 291108 40480
rect 291160 40468 291166 40520
rect 300854 40468 300860 40520
rect 300912 40508 300918 40520
rect 302142 40508 302148 40520
rect 300912 40480 302148 40508
rect 300912 40468 300918 40480
rect 302142 40468 302148 40480
rect 302200 40468 302206 40520
rect 283006 40332 283012 40384
rect 283064 40372 283070 40384
rect 284202 40372 284208 40384
rect 283064 40344 284208 40372
rect 283064 40332 283070 40344
rect 284202 40332 284208 40344
rect 284260 40332 284266 40384
rect 309137 40375 309195 40381
rect 309137 40341 309149 40375
rect 309183 40372 309195 40375
rect 313458 40372 313464 40384
rect 309183 40344 313464 40372
rect 309183 40341 309195 40344
rect 309137 40335 309195 40341
rect 313458 40332 313464 40344
rect 313516 40332 313522 40384
rect 335446 40332 335452 40384
rect 335504 40372 335510 40384
rect 336642 40372 336648 40384
rect 335504 40344 336648 40372
rect 335504 40332 335510 40344
rect 336642 40332 336648 40344
rect 336700 40332 336706 40384
rect 64874 40128 64880 40180
rect 64932 40168 64938 40180
rect 66162 40168 66168 40180
rect 64932 40140 66168 40168
rect 64932 40128 64938 40140
rect 66162 40128 66168 40140
rect 66220 40128 66226 40180
rect 66070 40060 66076 40112
rect 66128 40100 66134 40112
rect 66898 40100 66904 40112
rect 66128 40072 66904 40100
rect 66128 40060 66134 40072
rect 66898 40060 66904 40072
rect 66956 40060 66962 40112
rect 70854 40060 70860 40112
rect 70912 40100 70918 40112
rect 71682 40100 71688 40112
rect 70912 40072 71688 40100
rect 70912 40060 70918 40072
rect 71682 40060 71688 40072
rect 71740 40060 71746 40112
rect 72050 40060 72056 40112
rect 72108 40100 72114 40112
rect 73062 40100 73068 40112
rect 72108 40072 73068 40100
rect 72108 40060 72114 40072
rect 73062 40060 73068 40072
rect 73120 40060 73126 40112
rect 80422 40060 80428 40112
rect 80480 40100 80486 40112
rect 81342 40100 81348 40112
rect 80480 40072 81348 40100
rect 80480 40060 80486 40072
rect 81342 40060 81348 40072
rect 81400 40060 81406 40112
rect 82814 40060 82820 40112
rect 82872 40100 82878 40112
rect 84010 40100 84016 40112
rect 82872 40072 84016 40100
rect 82872 40060 82878 40072
rect 84010 40060 84016 40072
rect 84068 40060 84074 40112
rect 89898 40060 89904 40112
rect 89956 40100 89962 40112
rect 91002 40100 91008 40112
rect 89956 40072 91008 40100
rect 89956 40060 89962 40072
rect 91002 40060 91008 40072
rect 91060 40060 91066 40112
rect 91094 40060 91100 40112
rect 91152 40100 91158 40112
rect 92382 40100 92388 40112
rect 91152 40072 92388 40100
rect 91152 40060 91158 40072
rect 92382 40060 92388 40072
rect 92440 40060 92446 40112
rect 97074 40060 97080 40112
rect 97132 40100 97138 40112
rect 97902 40100 97908 40112
rect 97132 40072 97908 40100
rect 97132 40060 97138 40072
rect 97902 40060 97908 40072
rect 97960 40060 97966 40112
rect 98270 40060 98276 40112
rect 98328 40100 98334 40112
rect 99282 40100 99288 40112
rect 98328 40072 99288 40100
rect 98328 40060 98334 40072
rect 99282 40060 99288 40072
rect 99340 40060 99346 40112
rect 99466 40060 99472 40112
rect 99524 40100 99530 40112
rect 100662 40100 100668 40112
rect 99524 40072 100668 40100
rect 99524 40060 99530 40072
rect 100662 40060 100668 40072
rect 100720 40060 100726 40112
rect 105446 40060 105452 40112
rect 105504 40100 105510 40112
rect 106182 40100 106188 40112
rect 105504 40072 106188 40100
rect 105504 40060 105510 40072
rect 106182 40060 106188 40072
rect 106240 40060 106246 40112
rect 106642 40060 106648 40112
rect 106700 40100 106706 40112
rect 107562 40100 107568 40112
rect 106700 40072 107568 40100
rect 106700 40060 106706 40072
rect 107562 40060 107568 40072
rect 107620 40060 107626 40112
rect 107838 40060 107844 40112
rect 107896 40100 107902 40112
rect 108942 40100 108948 40112
rect 107896 40072 108948 40100
rect 107896 40060 107902 40072
rect 108942 40060 108948 40072
rect 109000 40060 109006 40112
rect 109034 40060 109040 40112
rect 109092 40100 109098 40112
rect 110322 40100 110328 40112
rect 109092 40072 110328 40100
rect 109092 40060 109098 40072
rect 110322 40060 110328 40072
rect 110380 40060 110386 40112
rect 113726 40060 113732 40112
rect 113784 40100 113790 40112
rect 114462 40100 114468 40112
rect 113784 40072 114468 40100
rect 113784 40060 113790 40072
rect 114462 40060 114468 40072
rect 114520 40060 114526 40112
rect 114922 40060 114928 40112
rect 114980 40100 114986 40112
rect 115842 40100 115848 40112
rect 114980 40072 115848 40100
rect 114980 40060 114986 40072
rect 115842 40060 115848 40072
rect 115900 40060 115906 40112
rect 116118 40060 116124 40112
rect 116176 40100 116182 40112
rect 117222 40100 117228 40112
rect 116176 40072 117228 40100
rect 116176 40060 116182 40072
rect 117222 40060 117228 40072
rect 117280 40060 117286 40112
rect 117314 40060 117320 40112
rect 117372 40100 117378 40112
rect 118602 40100 118608 40112
rect 117372 40072 118608 40100
rect 117372 40060 117378 40072
rect 118602 40060 118608 40072
rect 118660 40060 118666 40112
rect 124490 40060 124496 40112
rect 124548 40100 124554 40112
rect 125502 40100 125508 40112
rect 124548 40072 125508 40100
rect 124548 40060 124554 40072
rect 125502 40060 125508 40072
rect 125560 40060 125566 40112
rect 125686 40060 125692 40112
rect 125744 40100 125750 40112
rect 126790 40100 126796 40112
rect 125744 40072 126796 40100
rect 125744 40060 125750 40072
rect 126790 40060 126796 40072
rect 126848 40060 126854 40112
rect 132862 40060 132868 40112
rect 132920 40100 132926 40112
rect 133782 40100 133788 40112
rect 132920 40072 133788 40100
rect 132920 40060 132926 40072
rect 133782 40060 133788 40072
rect 133840 40060 133846 40112
rect 134058 40060 134064 40112
rect 134116 40100 134122 40112
rect 135162 40100 135168 40112
rect 134116 40072 135168 40100
rect 134116 40060 134122 40072
rect 135162 40060 135168 40072
rect 135220 40060 135226 40112
rect 135254 40060 135260 40112
rect 135312 40100 135318 40112
rect 136542 40100 136548 40112
rect 135312 40072 136548 40100
rect 135312 40060 135318 40072
rect 136542 40060 136548 40072
rect 136600 40060 136606 40112
rect 141142 40060 141148 40112
rect 141200 40100 141206 40112
rect 142062 40100 142068 40112
rect 141200 40072 142068 40100
rect 141200 40060 141206 40072
rect 142062 40060 142068 40072
rect 142120 40060 142126 40112
rect 142338 40060 142344 40112
rect 142396 40100 142402 40112
rect 143442 40100 143448 40112
rect 142396 40072 143448 40100
rect 142396 40060 142402 40072
rect 143442 40060 143448 40072
rect 143500 40060 143506 40112
rect 143534 40060 143540 40112
rect 143592 40100 143598 40112
rect 144822 40100 144828 40112
rect 143592 40072 144828 40100
rect 143592 40060 143598 40072
rect 144822 40060 144828 40072
rect 144880 40060 144886 40112
rect 149514 40060 149520 40112
rect 149572 40100 149578 40112
rect 150342 40100 150348 40112
rect 149572 40072 150348 40100
rect 149572 40060 149578 40072
rect 150342 40060 150348 40072
rect 150400 40060 150406 40112
rect 150710 40060 150716 40112
rect 150768 40100 150774 40112
rect 151722 40100 151728 40112
rect 150768 40072 151728 40100
rect 150768 40060 150774 40072
rect 151722 40060 151728 40072
rect 151780 40060 151786 40112
rect 157886 40060 157892 40112
rect 157944 40100 157950 40112
rect 158622 40100 158628 40112
rect 157944 40072 158628 40100
rect 157944 40060 157950 40072
rect 158622 40060 158628 40072
rect 158680 40060 158686 40112
rect 160278 40060 160284 40112
rect 160336 40100 160342 40112
rect 161382 40100 161388 40112
rect 160336 40072 161388 40100
rect 160336 40060 160342 40072
rect 161382 40060 161388 40072
rect 161440 40060 161446 40112
rect 161474 40060 161480 40112
rect 161532 40100 161538 40112
rect 162762 40100 162768 40112
rect 161532 40072 162768 40100
rect 161532 40060 161538 40072
rect 162762 40060 162768 40072
rect 162820 40060 162826 40112
rect 166166 40060 166172 40112
rect 166224 40100 166230 40112
rect 166902 40100 166908 40112
rect 166224 40072 166908 40100
rect 166224 40060 166230 40072
rect 166902 40060 166908 40072
rect 166960 40060 166966 40112
rect 168558 40060 168564 40112
rect 168616 40100 168622 40112
rect 169662 40100 169668 40112
rect 168616 40072 169668 40100
rect 168616 40060 168622 40072
rect 169662 40060 169668 40072
rect 169720 40060 169726 40112
rect 169754 40060 169760 40112
rect 169812 40100 169818 40112
rect 170950 40100 170956 40112
rect 169812 40072 170956 40100
rect 169812 40060 169818 40072
rect 170950 40060 170956 40072
rect 171008 40060 171014 40112
rect 175734 40060 175740 40112
rect 175792 40100 175798 40112
rect 176562 40100 176568 40112
rect 175792 40072 176568 40100
rect 175792 40060 175798 40072
rect 176562 40060 176568 40072
rect 176620 40060 176626 40112
rect 176930 40060 176936 40112
rect 176988 40100 176994 40112
rect 177942 40100 177948 40112
rect 176988 40072 177948 40100
rect 176988 40060 176994 40072
rect 177942 40060 177948 40072
rect 178000 40060 178006 40112
rect 178126 40060 178132 40112
rect 178184 40100 178190 40112
rect 179322 40100 179328 40112
rect 178184 40072 179328 40100
rect 178184 40060 178190 40072
rect 179322 40060 179328 40072
rect 179380 40060 179386 40112
rect 185302 40060 185308 40112
rect 185360 40100 185366 40112
rect 186222 40100 186228 40112
rect 185360 40072 186228 40100
rect 185360 40060 185366 40072
rect 186222 40060 186228 40072
rect 186280 40060 186286 40112
rect 186498 40060 186504 40112
rect 186556 40100 186562 40112
rect 187602 40100 187608 40112
rect 186556 40072 187608 40100
rect 186556 40060 186562 40072
rect 187602 40060 187608 40072
rect 187660 40060 187666 40112
rect 193582 40060 193588 40112
rect 193640 40100 193646 40112
rect 194502 40100 194508 40112
rect 193640 40072 194508 40100
rect 193640 40060 193646 40072
rect 194502 40060 194508 40072
rect 194560 40060 194566 40112
rect 195974 40060 195980 40112
rect 196032 40100 196038 40112
rect 197262 40100 197268 40112
rect 196032 40072 197268 40100
rect 196032 40060 196038 40072
rect 197262 40060 197268 40072
rect 197320 40060 197326 40112
rect 201954 40060 201960 40112
rect 202012 40100 202018 40112
rect 202782 40100 202788 40112
rect 202012 40072 202788 40100
rect 202012 40060 202018 40072
rect 202782 40060 202788 40072
rect 202840 40060 202846 40112
rect 203150 40060 203156 40112
rect 203208 40100 203214 40112
rect 204162 40100 204168 40112
rect 203208 40072 204168 40100
rect 203208 40060 203214 40072
rect 204162 40060 204168 40072
rect 204220 40060 204226 40112
rect 204346 40060 204352 40112
rect 204404 40100 204410 40112
rect 205542 40100 205548 40112
rect 204404 40072 205548 40100
rect 204404 40060 204410 40072
rect 205542 40060 205548 40072
rect 205600 40060 205606 40112
rect 211522 40060 211528 40112
rect 211580 40100 211586 40112
rect 212442 40100 212448 40112
rect 211580 40072 212448 40100
rect 211580 40060 211586 40072
rect 212442 40060 212448 40072
rect 212500 40060 212506 40112
rect 212718 40060 212724 40112
rect 212776 40100 212782 40112
rect 213822 40100 213828 40112
rect 212776 40072 213828 40100
rect 212776 40060 212782 40072
rect 213822 40060 213828 40072
rect 213880 40060 213886 40112
rect 213914 40060 213920 40112
rect 213972 40100 213978 40112
rect 215202 40100 215208 40112
rect 213972 40072 215208 40100
rect 213972 40060 213978 40072
rect 215202 40060 215208 40072
rect 215260 40060 215266 40112
rect 218606 40060 218612 40112
rect 218664 40100 218670 40112
rect 219342 40100 219348 40112
rect 218664 40072 219348 40100
rect 218664 40060 218670 40072
rect 219342 40060 219348 40072
rect 219400 40060 219406 40112
rect 220998 40060 221004 40112
rect 221056 40100 221062 40112
rect 222102 40100 222108 40112
rect 221056 40072 222108 40100
rect 221056 40060 221062 40072
rect 222102 40060 222108 40072
rect 222160 40060 222166 40112
rect 222194 40060 222200 40112
rect 222252 40100 222258 40112
rect 223482 40100 223488 40112
rect 222252 40072 223488 40100
rect 222252 40060 222258 40072
rect 223482 40060 223488 40072
rect 223540 40060 223546 40112
rect 228174 40060 228180 40112
rect 228232 40100 228238 40112
rect 229002 40100 229008 40112
rect 228232 40072 229008 40100
rect 228232 40060 228238 40072
rect 229002 40060 229008 40072
rect 229060 40060 229066 40112
rect 229370 40060 229376 40112
rect 229428 40100 229434 40112
rect 230382 40100 230388 40112
rect 229428 40072 230388 40100
rect 229428 40060 229434 40072
rect 230382 40060 230388 40072
rect 230440 40060 230446 40112
rect 230566 40060 230572 40112
rect 230624 40100 230630 40112
rect 231670 40100 231676 40112
rect 230624 40072 231676 40100
rect 230624 40060 230630 40072
rect 231670 40060 231676 40072
rect 231728 40060 231734 40112
rect 237742 40060 237748 40112
rect 237800 40100 237806 40112
rect 238662 40100 238668 40112
rect 237800 40072 238668 40100
rect 237800 40060 237806 40072
rect 238662 40060 238668 40072
rect 238720 40060 238726 40112
rect 238938 40060 238944 40112
rect 238996 40100 239002 40112
rect 240042 40100 240048 40112
rect 238996 40072 240048 40100
rect 238996 40060 239002 40072
rect 240042 40060 240048 40072
rect 240100 40060 240106 40112
rect 240134 40060 240140 40112
rect 240192 40100 240198 40112
rect 241422 40100 241428 40112
rect 240192 40072 241428 40100
rect 240192 40060 240198 40072
rect 241422 40060 241428 40072
rect 241480 40060 241486 40112
rect 246022 40060 246028 40112
rect 246080 40100 246086 40112
rect 246942 40100 246948 40112
rect 246080 40072 246948 40100
rect 246080 40060 246086 40072
rect 246942 40060 246948 40072
rect 247000 40060 247006 40112
rect 254394 40060 254400 40112
rect 254452 40100 254458 40112
rect 255222 40100 255228 40112
rect 254452 40072 255228 40100
rect 254452 40060 254458 40072
rect 255222 40060 255228 40072
rect 255280 40060 255286 40112
rect 255590 40060 255596 40112
rect 255648 40100 255654 40112
rect 256602 40100 256608 40112
rect 255648 40072 256608 40100
rect 255648 40060 255654 40072
rect 256602 40060 256608 40072
rect 256660 40060 256666 40112
rect 256786 40060 256792 40112
rect 256844 40100 256850 40112
rect 257982 40100 257988 40112
rect 256844 40072 257988 40100
rect 256844 40060 256850 40072
rect 257982 40060 257988 40072
rect 258040 40060 258046 40112
rect 262766 40060 262772 40112
rect 262824 40100 262830 40112
rect 263502 40100 263508 40112
rect 262824 40072 263508 40100
rect 262824 40060 262830 40072
rect 263502 40060 263508 40072
rect 263560 40060 263566 40112
rect 263962 40060 263968 40112
rect 264020 40100 264026 40112
rect 264882 40100 264888 40112
rect 264020 40072 264888 40100
rect 264020 40060 264026 40072
rect 264882 40060 264888 40072
rect 264940 40060 264946 40112
rect 265158 40060 265164 40112
rect 265216 40100 265222 40112
rect 266262 40100 266268 40112
rect 265216 40072 266268 40100
rect 265216 40060 265222 40072
rect 266262 40060 266268 40072
rect 266320 40060 266326 40112
rect 271046 40060 271052 40112
rect 271104 40100 271110 40112
rect 272518 40100 272524 40112
rect 271104 40072 272524 40100
rect 271104 40060 271110 40072
rect 272518 40060 272524 40072
rect 272576 40060 272582 40112
rect 274634 40060 274640 40112
rect 274692 40100 274698 40112
rect 275830 40100 275836 40112
rect 274692 40072 275836 40100
rect 274692 40060 274698 40072
rect 275830 40060 275836 40072
rect 275888 40060 275894 40112
rect 281810 40060 281816 40112
rect 281868 40100 281874 40112
rect 282822 40100 282828 40112
rect 281868 40072 282828 40100
rect 281868 40060 281874 40072
rect 282822 40060 282828 40072
rect 282880 40060 282886 40112
rect 291378 40060 291384 40112
rect 291436 40100 291442 40112
rect 292482 40100 292488 40112
rect 291436 40072 292488 40100
rect 291436 40060 291442 40072
rect 292482 40060 292488 40072
rect 292540 40060 292546 40112
rect 292574 40060 292580 40112
rect 292632 40100 292638 40112
rect 293862 40100 293868 40112
rect 292632 40072 293868 40100
rect 292632 40060 292638 40072
rect 293862 40060 293868 40072
rect 293920 40060 293926 40112
rect 306834 40060 306840 40112
rect 306892 40100 306898 40112
rect 307662 40100 307668 40112
rect 306892 40072 307668 40100
rect 306892 40060 306898 40072
rect 307662 40060 307668 40072
rect 307720 40060 307726 40112
rect 308030 40060 308036 40112
rect 308088 40100 308094 40112
rect 309042 40100 309048 40112
rect 308088 40072 309048 40100
rect 308088 40060 308094 40072
rect 309042 40060 309048 40072
rect 309100 40060 309106 40112
rect 309226 40060 309232 40112
rect 309284 40100 309290 40112
rect 311158 40100 311164 40112
rect 309284 40072 311164 40100
rect 309284 40060 309290 40072
rect 311158 40060 311164 40072
rect 311216 40060 311222 40112
rect 315206 40060 315212 40112
rect 315264 40100 315270 40112
rect 315942 40100 315948 40112
rect 315264 40072 315948 40100
rect 315264 40060 315270 40072
rect 315942 40060 315948 40072
rect 316000 40060 316006 40112
rect 317598 40060 317604 40112
rect 317656 40100 317662 40112
rect 318702 40100 318708 40112
rect 317656 40072 318708 40100
rect 317656 40060 317662 40072
rect 318702 40060 318708 40072
rect 318760 40060 318766 40112
rect 323486 40060 323492 40112
rect 323544 40100 323550 40112
rect 324222 40100 324228 40112
rect 323544 40072 324228 40100
rect 323544 40060 323550 40072
rect 324222 40060 324228 40072
rect 324280 40060 324286 40112
rect 325878 40060 325884 40112
rect 325936 40100 325942 40112
rect 326982 40100 326988 40112
rect 325936 40072 326988 40100
rect 325936 40060 325942 40072
rect 326982 40060 326988 40072
rect 327040 40060 327046 40112
rect 342622 40060 342628 40112
rect 342680 40100 342686 40112
rect 343542 40100 343548 40112
rect 342680 40072 343548 40100
rect 342680 40060 342686 40072
rect 343542 40060 343548 40072
rect 343600 40060 343606 40112
rect 350902 40060 350908 40112
rect 350960 40100 350966 40112
rect 351822 40100 351828 40112
rect 350960 40072 351828 40100
rect 350960 40060 350966 40072
rect 351822 40060 351828 40072
rect 351880 40060 351886 40112
rect 352098 40060 352104 40112
rect 352156 40100 352162 40112
rect 353202 40100 353208 40112
rect 352156 40072 353208 40100
rect 352156 40060 352162 40072
rect 353202 40060 353208 40072
rect 353260 40060 353266 40112
rect 353294 40060 353300 40112
rect 353352 40100 353358 40112
rect 354582 40100 354588 40112
rect 353352 40072 354588 40100
rect 353352 40060 353358 40072
rect 354582 40060 354588 40072
rect 354640 40060 354646 40112
rect 360470 40060 360476 40112
rect 360528 40100 360534 40112
rect 361482 40100 361488 40112
rect 360528 40072 361488 40100
rect 360528 40060 360534 40072
rect 361482 40060 361488 40072
rect 361540 40060 361546 40112
rect 361666 40060 361672 40112
rect 361724 40100 361730 40112
rect 362862 40100 362868 40112
rect 361724 40072 362868 40100
rect 361724 40060 361730 40072
rect 362862 40060 362868 40072
rect 362920 40060 362926 40112
rect 368842 40060 368848 40112
rect 368900 40100 368906 40112
rect 369762 40100 369768 40112
rect 368900 40072 369768 40100
rect 368900 40060 368906 40072
rect 369762 40060 369768 40072
rect 369820 40060 369826 40112
rect 375926 40060 375932 40112
rect 375984 40100 375990 40112
rect 376662 40100 376668 40112
rect 375984 40072 376668 40100
rect 375984 40060 375990 40072
rect 376662 40060 376668 40072
rect 376720 40060 376726 40112
rect 377122 40060 377128 40112
rect 377180 40100 377186 40112
rect 378042 40100 378048 40112
rect 377180 40072 378048 40100
rect 377180 40060 377186 40072
rect 378042 40060 378048 40072
rect 378100 40060 378106 40112
rect 379514 40060 379520 40112
rect 379572 40100 379578 40112
rect 380802 40100 380808 40112
rect 379572 40072 380808 40100
rect 379572 40060 379578 40072
rect 380802 40060 380808 40072
rect 380860 40060 380866 40112
rect 385494 40060 385500 40112
rect 385552 40100 385558 40112
rect 386322 40100 386328 40112
rect 385552 40072 386328 40100
rect 385552 40060 385558 40072
rect 386322 40060 386328 40072
rect 386380 40060 386386 40112
rect 386690 40060 386696 40112
rect 386748 40100 386754 40112
rect 387702 40100 387708 40112
rect 386748 40072 387708 40100
rect 386748 40060 386754 40072
rect 387702 40060 387708 40072
rect 387760 40060 387766 40112
rect 387886 40060 387892 40112
rect 387944 40100 387950 40112
rect 389082 40100 389088 40112
rect 387944 40072 389088 40100
rect 387944 40060 387950 40072
rect 389082 40060 389088 40072
rect 389140 40060 389146 40112
rect 394970 40060 394976 40112
rect 395028 40100 395034 40112
rect 395982 40100 395988 40112
rect 395028 40072 395988 40100
rect 395028 40060 395034 40072
rect 395982 40060 395988 40072
rect 396040 40060 396046 40112
rect 404538 40060 404544 40112
rect 404596 40100 404602 40112
rect 405642 40100 405648 40112
rect 404596 40072 405648 40100
rect 404596 40060 404602 40072
rect 405642 40060 405648 40072
rect 405700 40060 405706 40112
rect 405734 40060 405740 40112
rect 405792 40100 405798 40112
rect 406930 40100 406936 40112
rect 405792 40072 406936 40100
rect 405792 40060 405798 40072
rect 406930 40060 406936 40072
rect 406988 40060 406994 40112
rect 411714 40060 411720 40112
rect 411772 40100 411778 40112
rect 412542 40100 412548 40112
rect 411772 40072 412548 40100
rect 411772 40060 411778 40072
rect 412542 40060 412548 40072
rect 412600 40060 412606 40112
rect 412910 40060 412916 40112
rect 412968 40100 412974 40112
rect 413922 40100 413928 40112
rect 412968 40072 413928 40100
rect 412968 40060 412974 40072
rect 413922 40060 413928 40072
rect 413980 40060 413986 40112
rect 414106 40060 414112 40112
rect 414164 40100 414170 40112
rect 415302 40100 415308 40112
rect 414164 40072 415308 40100
rect 414164 40060 414170 40072
rect 415302 40060 415308 40072
rect 415360 40060 415366 40112
rect 420086 40060 420092 40112
rect 420144 40100 420150 40112
rect 420822 40100 420828 40112
rect 420144 40072 420828 40100
rect 420144 40060 420150 40072
rect 420822 40060 420828 40072
rect 420880 40060 420886 40112
rect 421190 40060 421196 40112
rect 421248 40100 421254 40112
rect 422202 40100 422208 40112
rect 421248 40072 422208 40100
rect 421248 40060 421254 40072
rect 422202 40060 422208 40072
rect 422260 40060 422266 40112
rect 422386 40060 422392 40112
rect 422444 40100 422450 40112
rect 423582 40100 423588 40112
rect 422444 40072 423588 40100
rect 422444 40060 422450 40072
rect 423582 40060 423588 40072
rect 423640 40060 423646 40112
rect 428366 40060 428372 40112
rect 428424 40100 428430 40112
rect 429102 40100 429108 40112
rect 428424 40072 429108 40100
rect 428424 40060 428430 40072
rect 429102 40060 429108 40072
rect 429160 40060 429166 40112
rect 429562 40060 429568 40112
rect 429620 40100 429626 40112
rect 430482 40100 430488 40112
rect 429620 40072 430488 40100
rect 429620 40060 429626 40072
rect 430482 40060 430488 40072
rect 430540 40060 430546 40112
rect 430758 40060 430764 40112
rect 430816 40100 430822 40112
rect 431862 40100 431868 40112
rect 430816 40072 431868 40100
rect 430816 40060 430822 40072
rect 431862 40060 431868 40072
rect 431920 40060 431926 40112
rect 431954 40060 431960 40112
rect 432012 40100 432018 40112
rect 433150 40100 433156 40112
rect 432012 40072 433156 40100
rect 432012 40060 432018 40072
rect 433150 40060 433156 40072
rect 433208 40060 433214 40112
rect 437934 40060 437940 40112
rect 437992 40100 437998 40112
rect 438762 40100 438768 40112
rect 437992 40072 438768 40100
rect 437992 40060 437998 40072
rect 438762 40060 438768 40072
rect 438820 40060 438826 40112
rect 439130 40060 439136 40112
rect 439188 40100 439194 40112
rect 440142 40100 440148 40112
rect 439188 40072 440148 40100
rect 439188 40060 439194 40072
rect 440142 40060 440148 40072
rect 440200 40060 440206 40112
rect 440326 40060 440332 40112
rect 440384 40100 440390 40112
rect 441522 40100 441528 40112
rect 440384 40072 441528 40100
rect 440384 40060 440390 40072
rect 441522 40060 441528 40072
rect 441580 40060 441586 40112
rect 446214 40060 446220 40112
rect 446272 40100 446278 40112
rect 447042 40100 447048 40112
rect 446272 40072 447048 40100
rect 446272 40060 446278 40072
rect 447042 40060 447048 40072
rect 447100 40060 447106 40112
rect 447410 40060 447416 40112
rect 447468 40100 447474 40112
rect 448422 40100 448428 40112
rect 447468 40072 448428 40100
rect 447468 40060 447474 40072
rect 448422 40060 448428 40072
rect 448480 40060 448486 40112
rect 448606 40060 448612 40112
rect 448664 40100 448670 40112
rect 449710 40100 449716 40112
rect 448664 40072 449716 40100
rect 448664 40060 448670 40072
rect 449710 40060 449716 40072
rect 449768 40060 449774 40112
rect 455782 40060 455788 40112
rect 455840 40100 455846 40112
rect 456702 40100 456708 40112
rect 455840 40072 456708 40100
rect 455840 40060 455846 40072
rect 456702 40060 456708 40072
rect 456760 40060 456766 40112
rect 456978 40060 456984 40112
rect 457036 40100 457042 40112
rect 458082 40100 458088 40112
rect 457036 40072 458088 40100
rect 457036 40060 457042 40072
rect 458082 40060 458088 40072
rect 458140 40060 458146 40112
rect 458174 40060 458180 40112
rect 458232 40100 458238 40112
rect 459462 40100 459468 40112
rect 458232 40072 459468 40100
rect 458232 40060 458238 40072
rect 459462 40060 459468 40072
rect 459520 40060 459526 40112
rect 464154 40060 464160 40112
rect 464212 40100 464218 40112
rect 464982 40100 464988 40112
rect 464212 40072 464988 40100
rect 464212 40060 464218 40072
rect 464982 40060 464988 40072
rect 465040 40060 465046 40112
rect 465350 40060 465356 40112
rect 465408 40100 465414 40112
rect 466362 40100 466368 40112
rect 465408 40072 466368 40100
rect 465408 40060 465414 40072
rect 466362 40060 466368 40072
rect 466420 40060 466426 40112
rect 466546 40060 466552 40112
rect 466604 40100 466610 40112
rect 467742 40100 467748 40112
rect 466604 40072 467748 40100
rect 466604 40060 466610 40072
rect 467742 40060 467748 40072
rect 467800 40060 467806 40112
rect 472434 40060 472440 40112
rect 472492 40100 472498 40112
rect 473262 40100 473268 40112
rect 472492 40072 473268 40100
rect 472492 40060 472498 40072
rect 473262 40060 473268 40072
rect 473320 40060 473326 40112
rect 473630 40060 473636 40112
rect 473688 40100 473694 40112
rect 474642 40100 474648 40112
rect 473688 40072 474648 40100
rect 473688 40060 473694 40072
rect 474642 40060 474648 40072
rect 474700 40060 474706 40112
rect 480806 40060 480812 40112
rect 480864 40100 480870 40112
rect 481542 40100 481548 40112
rect 480864 40072 481548 40100
rect 480864 40060 480870 40072
rect 481542 40060 481548 40072
rect 481600 40060 481606 40112
rect 483198 40060 483204 40112
rect 483256 40100 483262 40112
rect 484302 40100 484308 40112
rect 483256 40072 484308 40100
rect 483256 40060 483262 40072
rect 484302 40060 484308 40072
rect 484360 40060 484366 40112
rect 484394 40060 484400 40112
rect 484452 40100 484458 40112
rect 485590 40100 485596 40112
rect 484452 40072 485596 40100
rect 484452 40060 484458 40072
rect 485590 40060 485596 40072
rect 485648 40060 485654 40112
rect 490374 40060 490380 40112
rect 490432 40100 490438 40112
rect 491202 40100 491208 40112
rect 490432 40072 491208 40100
rect 490432 40060 490438 40072
rect 491202 40060 491208 40072
rect 491260 40060 491266 40112
rect 491570 40060 491576 40112
rect 491628 40100 491634 40112
rect 492582 40100 492588 40112
rect 491628 40072 492588 40100
rect 491628 40060 491634 40072
rect 492582 40060 492588 40072
rect 492640 40060 492646 40112
rect 492766 40060 492772 40112
rect 492824 40100 492830 40112
rect 493962 40100 493968 40112
rect 492824 40072 493968 40100
rect 492824 40060 492830 40072
rect 493962 40060 493968 40072
rect 494020 40060 494026 40112
rect 498654 40060 498660 40112
rect 498712 40100 498718 40112
rect 499482 40100 499488 40112
rect 498712 40072 499488 40100
rect 498712 40060 498718 40072
rect 499482 40060 499488 40072
rect 499540 40060 499546 40112
rect 499850 40060 499856 40112
rect 499908 40100 499914 40112
rect 500862 40100 500868 40112
rect 499908 40072 500868 40100
rect 499908 40060 499914 40072
rect 500862 40060 500868 40072
rect 500920 40060 500926 40112
rect 508222 40060 508228 40112
rect 508280 40100 508286 40112
rect 509142 40100 509148 40112
rect 508280 40072 509148 40100
rect 508280 40060 508286 40072
rect 509142 40060 509148 40072
rect 509200 40060 509206 40112
rect 509418 40060 509424 40112
rect 509476 40100 509482 40112
rect 510522 40100 510528 40112
rect 509476 40072 510528 40100
rect 509476 40060 509482 40072
rect 510522 40060 510528 40072
rect 510580 40060 510586 40112
rect 510614 40060 510620 40112
rect 510672 40100 510678 40112
rect 511902 40100 511908 40112
rect 510672 40072 511908 40100
rect 510672 40060 510678 40072
rect 511902 40060 511908 40072
rect 511960 40060 511966 40112
rect 516594 40060 516600 40112
rect 516652 40100 516658 40112
rect 517422 40100 517428 40112
rect 516652 40072 517428 40100
rect 516652 40060 516658 40072
rect 517422 40060 517428 40072
rect 517480 40060 517486 40112
rect 517790 40060 517796 40112
rect 517848 40100 517854 40112
rect 518802 40100 518808 40112
rect 517848 40072 518808 40100
rect 517848 40060 517854 40072
rect 518802 40060 518808 40072
rect 518860 40060 518866 40112
rect 287790 39448 287796 39500
rect 287848 39488 287854 39500
rect 347774 39488 347780 39500
rect 287848 39460 347780 39488
rect 287848 39448 287854 39460
rect 347774 39448 347780 39460
rect 347832 39448 347838 39500
rect 73246 39380 73252 39432
rect 73304 39420 73310 39432
rect 133874 39420 133880 39432
rect 73304 39392 133880 39420
rect 73304 39380 73310 39392
rect 133874 39380 133880 39392
rect 133932 39380 133938 39432
rect 159082 39380 159088 39432
rect 159140 39420 159146 39432
rect 219434 39420 219440 39432
rect 159140 39392 219440 39420
rect 159140 39380 159146 39392
rect 219434 39380 219440 39392
rect 219492 39380 219498 39432
rect 226978 39380 226984 39432
rect 227036 39420 227042 39432
rect 287054 39420 287060 39432
rect 227036 39392 287060 39420
rect 227036 39380 227042 39392
rect 287054 39380 287060 39392
rect 287112 39380 287118 39432
rect 319898 39380 319904 39432
rect 319956 39420 319962 39432
rect 380894 39420 380900 39432
rect 319956 39392 380900 39420
rect 319956 39380 319962 39392
rect 380894 39380 380900 39392
rect 380952 39380 380958 39432
rect 126882 39312 126888 39364
rect 126940 39352 126946 39364
rect 187694 39352 187700 39364
rect 126940 39324 187700 39352
rect 126940 39312 126946 39324
rect 187694 39312 187700 39324
rect 187752 39312 187758 39364
rect 194778 39312 194784 39364
rect 194836 39352 194842 39364
rect 255314 39352 255320 39364
rect 194836 39324 255320 39352
rect 194836 39312 194842 39324
rect 255314 39312 255320 39324
rect 255372 39312 255378 39364
rect 259178 39312 259184 39364
rect 259236 39352 259242 39364
rect 320174 39352 320180 39364
rect 259236 39324 320180 39352
rect 259236 39312 259242 39324
rect 320174 39312 320180 39324
rect 320232 39312 320238 39364
rect 366450 39312 366456 39364
rect 366508 39352 366514 39364
rect 426434 39352 426440 39364
rect 366508 39324 426440 39352
rect 366508 39312 366514 39324
rect 426434 39312 426440 39324
rect 426492 39312 426498 39364
rect 433242 39312 433248 39364
rect 433300 39352 433306 39364
rect 494054 39352 494060 39364
rect 433300 39324 494060 39352
rect 433300 39312 433306 39324
rect 494054 39312 494060 39324
rect 494112 39312 494118 39364
rect 501046 39312 501052 39364
rect 501104 39352 501110 39364
rect 561674 39352 561680 39364
rect 501104 39324 561680 39352
rect 501104 39312 501110 39324
rect 561674 39312 561680 39324
rect 561732 39312 561738 39364
rect 434806 38604 434812 38616
rect 434767 38576 434812 38604
rect 434806 38564 434812 38576
rect 434864 38564 434870 38616
rect 187970 38020 187976 38072
rect 188028 38060 188034 38072
rect 248414 38060 248420 38072
rect 188028 38032 248420 38060
rect 188028 38020 188034 38032
rect 248414 38020 248420 38032
rect 248472 38020 248478 38072
rect 402146 38020 402152 38072
rect 402204 38060 402210 38072
rect 462314 38060 462320 38072
rect 402204 38032 462320 38060
rect 402204 38020 402210 38032
rect 462314 38020 462320 38032
rect 462372 38020 462378 38072
rect 123294 37952 123300 38004
rect 123352 37992 123358 38004
rect 183554 37992 183560 38004
rect 123352 37964 183560 37992
rect 123352 37952 123358 37964
rect 183554 37952 183560 37964
rect 183612 37952 183618 38004
rect 219802 37952 219808 38004
rect 219860 37992 219866 38004
rect 280154 37992 280160 38004
rect 219860 37964 280160 37992
rect 219860 37952 219866 37964
rect 280154 37952 280160 37964
rect 280212 37952 280218 38004
rect 280614 37952 280620 38004
rect 280672 37992 280678 38004
rect 340874 37992 340880 38004
rect 280672 37964 340880 37992
rect 280672 37952 280678 37964
rect 340874 37952 340880 37964
rect 340932 37952 340938 38004
rect 359274 37952 359280 38004
rect 359332 37992 359338 38004
rect 419534 37992 419540 38004
rect 359332 37964 419540 37992
rect 359332 37952 359338 37964
rect 419534 37952 419540 37964
rect 419592 37952 419598 38004
rect 76834 37884 76840 37936
rect 76892 37924 76898 37936
rect 138014 37924 138020 37936
rect 76892 37896 138020 37924
rect 76892 37884 76898 37896
rect 138014 37884 138020 37896
rect 138072 37884 138078 37936
rect 155494 37884 155500 37936
rect 155552 37924 155558 37936
rect 216674 37924 216680 37936
rect 155552 37896 216680 37924
rect 155552 37884 155558 37896
rect 216674 37884 216680 37896
rect 216732 37884 216738 37936
rect 248690 37884 248696 37936
rect 248748 37924 248754 37936
rect 309134 37924 309140 37936
rect 248748 37896 309140 37924
rect 248748 37884 248754 37896
rect 309134 37884 309140 37896
rect 309192 37884 309198 37936
rect 312814 37884 312820 37936
rect 312872 37924 312878 37936
rect 374086 37924 374092 37936
rect 312872 37896 374092 37924
rect 312872 37884 312878 37896
rect 374086 37884 374092 37896
rect 374144 37884 374150 37936
rect 450998 37884 451004 37936
rect 451056 37924 451062 37936
rect 511994 37924 512000 37936
rect 451056 37896 512000 37924
rect 451056 37884 451062 37896
rect 511994 37884 512000 37896
rect 512052 37884 512058 37936
rect 518986 37884 518992 37936
rect 519044 37924 519050 37936
rect 579614 37924 579620 37936
rect 519044 37896 579620 37924
rect 519044 37884 519050 37896
rect 579614 37884 579620 37896
rect 579672 37884 579678 37936
rect 184106 36660 184112 36712
rect 184164 36700 184170 36712
rect 244274 36700 244280 36712
rect 184164 36672 244280 36700
rect 184164 36660 184170 36672
rect 244274 36660 244280 36672
rect 244332 36660 244338 36712
rect 244826 36660 244832 36712
rect 244884 36700 244890 36712
rect 304994 36700 305000 36712
rect 244884 36672 305000 36700
rect 244884 36660 244890 36672
rect 304994 36660 305000 36672
rect 305052 36660 305058 36712
rect 305638 36660 305644 36712
rect 305696 36700 305702 36712
rect 365714 36700 365720 36712
rect 305696 36672 365720 36700
rect 305696 36660 305702 36672
rect 365714 36660 365720 36672
rect 365772 36660 365778 36712
rect 151906 36592 151912 36644
rect 151964 36632 151970 36644
rect 212534 36632 212540 36644
rect 151964 36604 212540 36632
rect 151964 36592 151970 36604
rect 212534 36592 212540 36604
rect 212592 36592 212598 36644
rect 277026 36592 277032 36644
rect 277084 36632 277090 36644
rect 338114 36632 338120 36644
rect 277084 36604 338120 36632
rect 277084 36592 277090 36604
rect 338114 36592 338120 36604
rect 338172 36592 338178 36644
rect 119706 36524 119712 36576
rect 119764 36564 119770 36576
rect 180794 36564 180800 36576
rect 119764 36536 180800 36564
rect 119764 36524 119770 36536
rect 180794 36524 180800 36536
rect 180852 36524 180858 36576
rect 216214 36524 216220 36576
rect 216272 36564 216278 36576
rect 277394 36564 277400 36576
rect 216272 36536 277400 36564
rect 216272 36524 216278 36536
rect 277394 36524 277400 36536
rect 277452 36524 277458 36576
rect 348510 36524 348516 36576
rect 348568 36564 348574 36576
rect 408494 36564 408500 36576
rect 348568 36536 408500 36564
rect 348568 36524 348574 36536
rect 408494 36524 408500 36536
rect 408552 36524 408558 36576
rect 415210 36524 415216 36576
rect 415268 36564 415274 36576
rect 476114 36564 476120 36576
rect 415268 36536 476120 36564
rect 415268 36524 415274 36536
rect 476114 36524 476120 36536
rect 476172 36524 476178 36576
rect 493870 36524 493876 36576
rect 493928 36564 493934 36576
rect 554774 36564 554780 36576
rect 493928 36536 554780 36564
rect 493928 36524 493934 36536
rect 554774 36524 554780 36536
rect 554832 36524 554838 36576
rect 213822 35300 213828 35352
rect 213880 35340 213886 35352
rect 273254 35340 273260 35352
rect 213880 35312 273260 35340
rect 213880 35300 213886 35312
rect 273254 35300 273260 35312
rect 273312 35300 273318 35352
rect 273438 35300 273444 35352
rect 273496 35340 273502 35352
rect 333974 35340 333980 35352
rect 273496 35312 333980 35340
rect 273496 35300 273502 35312
rect 333974 35300 333980 35312
rect 334032 35300 334038 35352
rect 117222 35232 117228 35284
rect 117280 35272 117286 35284
rect 176654 35272 176660 35284
rect 117280 35244 176660 35272
rect 117280 35232 117286 35244
rect 176654 35232 176660 35244
rect 176712 35232 176718 35284
rect 180702 35232 180708 35284
rect 180760 35272 180766 35284
rect 241514 35272 241520 35284
rect 180760 35244 241520 35272
rect 180760 35232 180766 35244
rect 241514 35232 241520 35244
rect 241572 35232 241578 35284
rect 302050 35232 302056 35284
rect 302108 35272 302114 35284
rect 362954 35272 362960 35284
rect 302108 35244 362960 35272
rect 302108 35232 302114 35244
rect 362954 35232 362960 35244
rect 363012 35232 363018 35284
rect 391842 35232 391848 35284
rect 391900 35272 391906 35284
rect 451274 35272 451280 35284
rect 391900 35244 451280 35272
rect 391900 35232 391906 35244
rect 451274 35232 451280 35244
rect 451332 35232 451338 35284
rect 148962 35164 148968 35216
rect 149020 35204 149026 35216
rect 209866 35204 209872 35216
rect 149020 35176 209872 35204
rect 149020 35164 149026 35176
rect 209866 35164 209872 35176
rect 209924 35164 209930 35216
rect 241330 35164 241336 35216
rect 241388 35204 241394 35216
rect 302234 35204 302240 35216
rect 241388 35176 302240 35204
rect 241388 35164 241394 35176
rect 302234 35164 302240 35176
rect 302292 35164 302298 35216
rect 342162 35164 342168 35216
rect 342220 35204 342226 35216
rect 401594 35204 401600 35216
rect 342220 35176 401600 35204
rect 342220 35164 342226 35176
rect 401594 35164 401600 35176
rect 401652 35164 401658 35216
rect 413922 35164 413928 35216
rect 413980 35204 413986 35216
rect 473354 35204 473360 35216
rect 413980 35176 473360 35204
rect 413980 35164 413986 35176
rect 473354 35164 473360 35176
rect 473412 35164 473418 35216
rect 511810 35164 511816 35216
rect 511868 35204 511874 35216
rect 571426 35204 571432 35216
rect 511868 35176 571432 35204
rect 511868 35164 511874 35176
rect 571426 35164 571432 35176
rect 571484 35164 571490 35216
rect 177942 33872 177948 33924
rect 178000 33912 178006 33924
rect 237374 33912 237380 33924
rect 178000 33884 237380 33912
rect 178000 33872 178006 33884
rect 237374 33872 237380 33884
rect 237432 33872 237438 33924
rect 238662 33872 238668 33924
rect 238720 33912 238726 33924
rect 298094 33912 298100 33924
rect 238720 33884 298100 33912
rect 238720 33872 238726 33884
rect 298094 33872 298100 33884
rect 298152 33872 298158 33924
rect 113082 33804 113088 33856
rect 113140 33844 113146 33856
rect 173894 33844 173900 33856
rect 113140 33816 173900 33844
rect 113140 33804 113146 33816
rect 173894 33804 173900 33816
rect 173952 33804 173958 33856
rect 205450 33804 205456 33856
rect 205508 33844 205514 33856
rect 266354 33844 266360 33856
rect 205508 33816 266360 33844
rect 205508 33804 205514 33816
rect 266354 33804 266360 33816
rect 266412 33804 266418 33856
rect 298462 33804 298468 33856
rect 298520 33844 298526 33856
rect 358814 33844 358820 33856
rect 298520 33816 358820 33844
rect 298520 33804 298526 33816
rect 358814 33804 358820 33816
rect 358872 33804 358878 33856
rect 383102 33804 383108 33856
rect 383160 33844 383166 33856
rect 383562 33844 383568 33856
rect 383160 33816 383568 33844
rect 383160 33804 383166 33816
rect 383562 33804 383568 33816
rect 383620 33804 383626 33856
rect 384942 33804 384948 33856
rect 385000 33844 385006 33856
rect 444374 33844 444380 33856
rect 385000 33816 444380 33844
rect 385000 33804 385006 33816
rect 444374 33804 444380 33816
rect 444432 33804 444438 33856
rect 449710 33804 449716 33856
rect 449768 33844 449774 33856
rect 509234 33844 509240 33856
rect 449768 33816 509240 33844
rect 449768 33804 449774 33816
rect 509234 33804 509240 33816
rect 509292 33804 509298 33856
rect 144730 33736 144736 33788
rect 144788 33776 144794 33788
rect 205634 33776 205640 33788
rect 144788 33748 205640 33776
rect 144788 33736 144794 33748
rect 205634 33736 205640 33748
rect 205692 33736 205698 33788
rect 270402 33736 270408 33788
rect 270460 33776 270466 33788
rect 331214 33776 331220 33788
rect 270460 33748 331220 33776
rect 270460 33736 270466 33748
rect 331214 33736 331220 33748
rect 331272 33736 331278 33788
rect 338022 33736 338028 33788
rect 338080 33776 338086 33788
rect 398926 33776 398932 33788
rect 338080 33748 398932 33776
rect 338080 33736 338086 33748
rect 398926 33736 398932 33748
rect 398984 33736 398990 33788
rect 502150 33736 502156 33788
rect 502208 33776 502214 33788
rect 563146 33776 563152 33788
rect 502208 33748 563152 33776
rect 502208 33736 502214 33748
rect 563146 33736 563152 33748
rect 563204 33736 563210 33788
rect 266538 32512 266544 32564
rect 266596 32552 266602 32564
rect 327074 32552 327080 32564
rect 266596 32524 327080 32552
rect 266596 32512 266602 32524
rect 327074 32512 327080 32524
rect 327132 32512 327138 32564
rect 142062 32444 142068 32496
rect 142120 32484 142126 32496
rect 201494 32484 201500 32496
rect 142120 32456 201500 32484
rect 142120 32444 142126 32456
rect 201494 32444 201500 32456
rect 201552 32444 201558 32496
rect 202782 32444 202788 32496
rect 202840 32484 202846 32496
rect 262214 32484 262220 32496
rect 202840 32456 262220 32484
rect 202840 32444 202846 32456
rect 262214 32444 262220 32456
rect 262272 32444 262278 32496
rect 295242 32444 295248 32496
rect 295300 32484 295306 32496
rect 356146 32484 356152 32496
rect 295300 32456 356152 32484
rect 295300 32444 295306 32456
rect 356146 32444 356152 32456
rect 356204 32444 356210 32496
rect 373902 32444 373908 32496
rect 373960 32484 373966 32496
rect 433334 32484 433340 32496
rect 373960 32456 433340 32484
rect 373960 32444 373966 32456
rect 433334 32444 433340 32456
rect 433392 32444 433398 32496
rect 445662 32444 445668 32496
rect 445720 32484 445726 32496
rect 505094 32484 505100 32496
rect 445720 32456 505100 32484
rect 445720 32444 445726 32456
rect 505094 32444 505100 32456
rect 505152 32444 505158 32496
rect 110322 32376 110328 32428
rect 110380 32416 110386 32428
rect 169754 32416 169760 32428
rect 110380 32388 169760 32416
rect 110380 32376 110386 32388
rect 169754 32376 169760 32388
rect 169812 32376 169818 32428
rect 170950 32376 170956 32428
rect 171008 32416 171014 32428
rect 230474 32416 230480 32428
rect 171008 32388 230480 32416
rect 171008 32376 171014 32388
rect 230474 32376 230480 32388
rect 230532 32376 230538 32428
rect 234522 32376 234528 32428
rect 234580 32416 234586 32428
rect 295334 32416 295340 32428
rect 234580 32388 295340 32416
rect 234580 32376 234586 32388
rect 295334 32376 295340 32388
rect 295392 32376 295398 32428
rect 327258 32376 327264 32428
rect 327316 32416 327322 32428
rect 387794 32416 387800 32428
rect 327316 32388 387800 32416
rect 327316 32376 327322 32388
rect 387794 32376 387800 32388
rect 387852 32376 387858 32428
rect 420822 32376 420828 32428
rect 420880 32416 420886 32428
rect 480254 32416 480260 32428
rect 420880 32388 480260 32416
rect 420880 32376 420886 32388
rect 480254 32376 480260 32388
rect 480312 32376 480318 32428
rect 495342 32376 495348 32428
rect 495400 32416 495406 32428
rect 554866 32416 554872 32428
rect 495400 32388 554872 32416
rect 495400 32376 495406 32388
rect 554866 32376 554872 32388
rect 554924 32376 554930 32428
rect 135162 31152 135168 31204
rect 135220 31192 135226 31204
rect 194594 31192 194600 31204
rect 135220 31164 194600 31192
rect 135220 31152 135226 31164
rect 194594 31152 194600 31164
rect 194652 31152 194658 31204
rect 106182 31084 106188 31136
rect 106240 31124 106246 31136
rect 167086 31124 167092 31136
rect 106240 31096 167092 31124
rect 106240 31084 106246 31096
rect 167086 31084 167092 31096
rect 167144 31084 167150 31136
rect 198642 31084 198648 31136
rect 198700 31124 198706 31136
rect 259454 31124 259460 31136
rect 198700 31096 259460 31124
rect 198700 31084 198706 31096
rect 259454 31084 259460 31096
rect 259512 31084 259518 31136
rect 263502 31084 263508 31136
rect 263560 31124 263566 31136
rect 322934 31124 322940 31136
rect 263560 31096 322940 31124
rect 263560 31084 263566 31096
rect 322934 31084 322940 31096
rect 322992 31084 322998 31136
rect 324222 31084 324228 31136
rect 324280 31124 324286 31136
rect 383654 31124 383660 31136
rect 324280 31096 383660 31124
rect 324280 31084 324286 31096
rect 383654 31084 383660 31096
rect 383712 31084 383718 31136
rect 492582 31084 492588 31136
rect 492640 31124 492646 31136
rect 552014 31124 552020 31136
rect 492640 31096 552020 31124
rect 492640 31084 492646 31096
rect 552014 31084 552020 31096
rect 552072 31084 552078 31136
rect 166902 31016 166908 31068
rect 166960 31056 166966 31068
rect 227806 31056 227812 31068
rect 166960 31028 227812 31056
rect 166960 31016 166966 31028
rect 227806 31016 227812 31028
rect 227864 31016 227870 31068
rect 231670 31016 231676 31068
rect 231728 31056 231734 31068
rect 291194 31056 291200 31068
rect 231728 31028 291200 31056
rect 231728 31016 231734 31028
rect 291194 31016 291200 31028
rect 291252 31016 291258 31068
rect 292482 31016 292488 31068
rect 292540 31056 292546 31068
rect 351914 31056 351920 31068
rect 292540 31028 351920 31056
rect 292540 31016 292546 31028
rect 351914 31016 351920 31028
rect 351972 31016 351978 31068
rect 371050 31016 371056 31068
rect 371108 31056 371114 31068
rect 430574 31056 430580 31068
rect 371108 31028 430580 31056
rect 371108 31016 371114 31028
rect 430574 31016 430580 31028
rect 430632 31016 430638 31068
rect 441430 31016 441436 31068
rect 441488 31056 441494 31068
rect 502426 31056 502432 31068
rect 441488 31028 502432 31056
rect 441488 31016 441494 31028
rect 502426 31016 502432 31028
rect 502484 31016 502490 31068
rect 523862 30268 523868 30320
rect 523920 30308 523926 30320
rect 580166 30308 580172 30320
rect 523920 30280 580172 30308
rect 523920 30268 523926 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 191742 29792 191748 29844
rect 191800 29832 191806 29844
rect 252646 29832 252652 29844
rect 191800 29804 252652 29832
rect 191800 29792 191806 29804
rect 252646 29792 252652 29804
rect 252704 29792 252710 29844
rect 131022 29724 131028 29776
rect 131080 29764 131086 29776
rect 191834 29764 191840 29776
rect 131080 29736 191840 29764
rect 131080 29724 131086 29736
rect 191834 29724 191840 29736
rect 191892 29724 191898 29776
rect 256602 29724 256608 29776
rect 256660 29764 256666 29776
rect 316034 29764 316040 29776
rect 256660 29736 316040 29764
rect 256660 29724 256666 29736
rect 316034 29724 316040 29736
rect 316092 29724 316098 29776
rect 102042 29656 102048 29708
rect 102100 29696 102106 29708
rect 162854 29696 162860 29708
rect 102100 29668 162860 29696
rect 102100 29656 102106 29668
rect 162854 29656 162860 29668
rect 162912 29656 162918 29708
rect 223390 29656 223396 29708
rect 223448 29696 223454 29708
rect 284294 29696 284300 29708
rect 223448 29668 284300 29696
rect 223448 29656 223454 29668
rect 284294 29656 284300 29668
rect 284352 29656 284358 29708
rect 406930 29656 406936 29708
rect 406988 29696 406994 29708
rect 466454 29696 466460 29708
rect 406988 29668 466460 29696
rect 406988 29656 406994 29668
rect 466454 29656 466460 29668
rect 466512 29656 466518 29708
rect 162670 29588 162676 29640
rect 162728 29628 162734 29640
rect 223574 29628 223580 29640
rect 162728 29600 223580 29628
rect 162728 29588 162734 29600
rect 223574 29588 223580 29600
rect 223632 29588 223638 29640
rect 284110 29588 284116 29640
rect 284168 29628 284174 29640
rect 345014 29628 345020 29640
rect 284168 29600 345020 29628
rect 284168 29588 284174 29600
rect 345014 29588 345020 29600
rect 345072 29588 345078 29640
rect 354490 29588 354496 29640
rect 354548 29628 354554 29640
rect 415394 29628 415400 29640
rect 354548 29600 415400 29628
rect 354548 29588 354554 29600
rect 415394 29588 415400 29600
rect 415452 29588 415458 29640
rect 438762 29588 438768 29640
rect 438820 29628 438826 29640
rect 498194 29628 498200 29640
rect 438820 29600 498200 29628
rect 438820 29588 438826 29600
rect 498194 29588 498200 29600
rect 498252 29588 498258 29640
rect 434806 29016 434812 29028
rect 434767 28988 434812 29016
rect 434806 28976 434812 28988
rect 434864 28976 434870 29028
rect 383286 28908 383292 28960
rect 383344 28948 383350 28960
rect 383473 28951 383531 28957
rect 383473 28948 383485 28951
rect 383344 28920 383485 28948
rect 383344 28908 383350 28920
rect 383473 28917 383485 28920
rect 383519 28917 383531 28951
rect 383473 28911 383531 28917
rect 272518 28296 272524 28348
rect 272576 28336 272582 28348
rect 331306 28336 331312 28348
rect 272576 28308 331312 28336
rect 272576 28296 272582 28308
rect 331306 28296 331312 28308
rect 331364 28296 331370 28348
rect 378042 28296 378048 28348
rect 378100 28336 378106 28348
rect 437474 28336 437480 28348
rect 378100 28308 437480 28336
rect 378100 28296 378106 28308
rect 437474 28296 437480 28308
rect 437532 28296 437538 28348
rect 488442 28296 488448 28348
rect 488500 28336 488506 28348
rect 547874 28336 547880 28348
rect 488500 28308 547880 28336
rect 488500 28296 488506 28308
rect 547874 28296 547880 28308
rect 547932 28296 547938 28348
rect 97902 28228 97908 28280
rect 97960 28268 97966 28280
rect 158806 28268 158812 28280
rect 97960 28240 158812 28268
rect 97960 28228 97966 28240
rect 158806 28228 158812 28240
rect 158864 28228 158870 28280
rect 165522 28228 165528 28280
rect 165580 28268 165586 28280
rect 226334 28268 226340 28280
rect 165580 28240 226340 28268
rect 165580 28228 165586 28240
rect 226334 28228 226340 28240
rect 226392 28228 226398 28280
rect 244182 28228 244188 28280
rect 244240 28268 244246 28280
rect 305086 28268 305092 28280
rect 244240 28240 305092 28268
rect 244240 28228 244246 28240
rect 305086 28228 305092 28240
rect 305144 28228 305150 28280
rect 329742 28228 329748 28280
rect 329800 28268 329806 28280
rect 390554 28268 390560 28280
rect 329800 28240 390560 28268
rect 329800 28228 329806 28240
rect 390554 28228 390560 28240
rect 390612 28228 390618 28280
rect 434622 28228 434628 28280
rect 434680 28268 434686 28280
rect 494146 28268 494152 28280
rect 434680 28240 494152 28268
rect 434680 28228 434686 28240
rect 494146 28228 494152 28240
rect 494204 28228 494210 28280
rect 398834 27548 398840 27600
rect 398892 27588 398898 27600
rect 398926 27588 398932 27600
rect 398892 27560 398932 27588
rect 398892 27548 398898 27560
rect 398926 27548 398932 27560
rect 398984 27548 398990 27600
rect 275830 26936 275836 26988
rect 275888 26976 275894 26988
rect 335354 26976 335360 26988
rect 275888 26948 335360 26976
rect 275888 26936 275894 26948
rect 335354 26936 335360 26948
rect 335412 26936 335418 26988
rect 353202 26936 353208 26988
rect 353260 26976 353266 26988
rect 412637 26979 412695 26985
rect 412637 26976 412649 26979
rect 353260 26948 412649 26976
rect 353260 26936 353266 26948
rect 412637 26945 412649 26948
rect 412683 26945 412695 26979
rect 412637 26939 412695 26945
rect 431862 26936 431868 26988
rect 431920 26976 431926 26988
rect 491294 26976 491300 26988
rect 431920 26948 491300 26976
rect 431920 26936 431926 26948
rect 491294 26936 491300 26948
rect 491352 26936 491358 26988
rect 93762 26868 93768 26920
rect 93820 26908 93826 26920
rect 154574 26908 154580 26920
rect 93820 26880 154580 26908
rect 93820 26868 93826 26880
rect 154574 26868 154580 26880
rect 154632 26868 154638 26920
rect 158622 26868 158628 26920
rect 158680 26908 158686 26920
rect 218146 26908 218152 26920
rect 158680 26880 218152 26908
rect 158680 26868 158686 26880
rect 218146 26868 218152 26880
rect 218204 26868 218210 26920
rect 237282 26868 237288 26920
rect 237340 26908 237346 26920
rect 296806 26908 296812 26920
rect 237340 26880 296812 26908
rect 237340 26868 237346 26880
rect 296806 26868 296812 26880
rect 296864 26868 296870 26920
rect 311802 26868 311808 26920
rect 311860 26908 311866 26920
rect 372706 26908 372712 26920
rect 311860 26880 372712 26908
rect 311860 26868 311866 26880
rect 372706 26868 372712 26880
rect 372764 26868 372770 26920
rect 409782 26868 409788 26920
rect 409840 26908 409846 26920
rect 469214 26908 469220 26920
rect 409840 26880 469220 26908
rect 409840 26868 409846 26880
rect 469214 26868 469220 26880
rect 469272 26868 469278 26920
rect 485590 26868 485596 26920
rect 485648 26908 485654 26920
rect 545114 26908 545120 26920
rect 485648 26880 545120 26908
rect 485648 26868 485654 26880
rect 545114 26868 545120 26880
rect 545172 26868 545178 26920
rect 317322 25576 317328 25628
rect 317380 25616 317386 25628
rect 376754 25616 376760 25628
rect 317380 25588 376760 25616
rect 317380 25576 317386 25588
rect 376754 25576 376760 25588
rect 376812 25576 376818 25628
rect 427722 25576 427728 25628
rect 427780 25616 427786 25628
rect 487154 25616 487160 25628
rect 427780 25588 487160 25616
rect 427780 25576 427786 25588
rect 487154 25576 487160 25588
rect 487212 25576 487218 25628
rect 91002 25508 91008 25560
rect 91060 25548 91066 25560
rect 150526 25548 150532 25560
rect 91060 25520 150532 25548
rect 91060 25508 91066 25520
rect 150526 25508 150532 25520
rect 150584 25508 150590 25560
rect 154482 25508 154488 25560
rect 154540 25548 154546 25560
rect 215294 25548 215300 25560
rect 154540 25520 215300 25548
rect 154540 25508 154546 25520
rect 215294 25508 215300 25520
rect 215352 25508 215358 25560
rect 226242 25508 226248 25560
rect 226300 25548 226306 25560
rect 287146 25548 287152 25560
rect 226300 25520 287152 25548
rect 226300 25508 226306 25520
rect 287146 25508 287152 25520
rect 287204 25508 287210 25560
rect 293770 25508 293776 25560
rect 293828 25548 293834 25560
rect 354674 25548 354680 25560
rect 293828 25520 354680 25548
rect 293828 25508 293834 25520
rect 354674 25508 354680 25520
rect 354732 25508 354738 25560
rect 362770 25508 362776 25560
rect 362828 25548 362834 25560
rect 423674 25548 423680 25560
rect 362828 25520 423680 25548
rect 362828 25508 362834 25520
rect 423674 25508 423680 25520
rect 423732 25508 423738 25560
rect 477402 25508 477408 25560
rect 477460 25548 477466 25560
rect 536834 25548 536840 25560
rect 477460 25520 536840 25548
rect 477460 25508 477466 25520
rect 536834 25508 536840 25520
rect 536892 25508 536898 25560
rect 285582 24148 285588 24200
rect 285640 24188 285646 24200
rect 346394 24188 346400 24200
rect 285640 24160 346400 24188
rect 285640 24148 285646 24160
rect 346394 24148 346400 24160
rect 346452 24148 346458 24200
rect 474642 24148 474648 24200
rect 474700 24188 474706 24200
rect 534074 24188 534080 24200
rect 474700 24160 534080 24188
rect 474700 24148 474706 24160
rect 534074 24148 534080 24160
rect 534132 24148 534138 24200
rect 86862 24080 86868 24132
rect 86920 24120 86926 24132
rect 147674 24120 147680 24132
rect 86920 24092 147680 24120
rect 86920 24080 86926 24092
rect 147674 24080 147680 24092
rect 147732 24080 147738 24132
rect 151722 24080 151728 24132
rect 151780 24120 151786 24132
rect 211154 24120 211160 24132
rect 151780 24092 211160 24120
rect 151780 24080 151786 24092
rect 211154 24080 211160 24092
rect 211212 24080 211218 24132
rect 212442 24080 212448 24132
rect 212500 24120 212506 24132
rect 271874 24120 271880 24132
rect 212500 24092 271880 24120
rect 212500 24080 212506 24092
rect 271874 24080 271880 24092
rect 271932 24080 271938 24132
rect 275922 24080 275928 24132
rect 275980 24120 275986 24132
rect 336734 24120 336740 24132
rect 275980 24092 336740 24120
rect 275980 24080 275986 24092
rect 336734 24080 336740 24092
rect 336792 24080 336798 24132
rect 344830 24080 344836 24132
rect 344888 24120 344894 24132
rect 404354 24120 404360 24132
rect 344888 24092 404360 24120
rect 344888 24080 344894 24092
rect 404354 24080 404360 24092
rect 404412 24080 404418 24132
rect 423490 24080 423496 24132
rect 423548 24120 423554 24132
rect 484394 24120 484400 24132
rect 423548 24092 484400 24120
rect 423548 24080 423554 24092
rect 484394 24080 484400 24092
rect 484452 24080 484458 24132
rect 278682 22788 278688 22840
rect 278740 22828 278746 22840
rect 339494 22828 339500 22840
rect 278740 22800 339500 22828
rect 278740 22788 278746 22800
rect 339494 22788 339500 22800
rect 339552 22788 339558 22840
rect 467742 22788 467748 22840
rect 467800 22828 467806 22840
rect 527174 22828 527180 22840
rect 467800 22800 527180 22828
rect 467800 22788 467806 22800
rect 527174 22788 527180 22800
rect 527232 22788 527238 22840
rect 84010 22720 84016 22772
rect 84068 22760 84074 22772
rect 143534 22760 143540 22772
rect 84068 22732 143540 22760
rect 84068 22720 84074 22732
rect 143534 22720 143540 22732
rect 143592 22720 143598 22772
rect 147582 22720 147588 22772
rect 147640 22760 147646 22772
rect 208394 22760 208400 22772
rect 147640 22732 208400 22760
rect 147640 22720 147646 22732
rect 208394 22720 208400 22732
rect 208452 22720 208458 22772
rect 215110 22720 215116 22772
rect 215168 22760 215174 22772
rect 276014 22760 276020 22772
rect 215168 22732 276020 22760
rect 215168 22720 215174 22732
rect 276014 22720 276020 22732
rect 276072 22720 276078 22772
rect 286962 22720 286968 22772
rect 287020 22760 287026 22772
rect 347866 22760 347872 22772
rect 287020 22732 347872 22760
rect 287020 22720 287026 22732
rect 347866 22720 347872 22732
rect 347924 22720 347930 22772
rect 351822 22720 351828 22772
rect 351880 22760 351886 22772
rect 411254 22760 411260 22772
rect 351880 22732 411260 22760
rect 351880 22720 351886 22732
rect 411254 22720 411260 22732
rect 411312 22720 411318 22772
rect 412542 22720 412548 22772
rect 412600 22760 412606 22772
rect 471974 22760 471980 22772
rect 412600 22732 471980 22760
rect 412600 22720 412606 22732
rect 471974 22720 471980 22732
rect 472032 22720 472038 22772
rect 383470 22012 383476 22024
rect 383431 21984 383476 22012
rect 383470 21972 383476 21984
rect 383528 21972 383534 22024
rect 419442 21428 419448 21480
rect 419500 21468 419506 21480
rect 478874 21468 478880 21480
rect 419500 21440 478880 21468
rect 419500 21428 419506 21440
rect 478874 21428 478880 21440
rect 478932 21428 478938 21480
rect 79962 21360 79968 21412
rect 80020 21400 80026 21412
rect 140774 21400 140780 21412
rect 80020 21372 140780 21400
rect 80020 21360 80026 21372
rect 140774 21360 140780 21372
rect 140832 21360 140838 21412
rect 144822 21360 144828 21412
rect 144880 21400 144886 21412
rect 204254 21400 204260 21412
rect 144880 21372 204260 21400
rect 144880 21360 144886 21372
rect 204254 21360 204260 21372
rect 204312 21360 204318 21412
rect 205542 21360 205548 21412
rect 205600 21400 205606 21412
rect 264974 21400 264980 21412
rect 205600 21372 264980 21400
rect 205600 21360 205606 21372
rect 264974 21360 264980 21372
rect 265032 21360 265038 21412
rect 269022 21360 269028 21412
rect 269080 21400 269086 21412
rect 329834 21400 329840 21412
rect 269080 21372 329840 21400
rect 269080 21360 269086 21372
rect 329834 21360 329840 21372
rect 329892 21360 329898 21412
rect 336550 21360 336556 21412
rect 336608 21400 336614 21412
rect 397454 21400 397460 21412
rect 336608 21372 397460 21400
rect 336608 21360 336614 21372
rect 397454 21360 397460 21372
rect 397512 21360 397518 21412
rect 470502 21360 470508 21412
rect 470560 21400 470566 21412
rect 529934 21400 529940 21412
rect 470560 21372 529940 21400
rect 470560 21360 470566 21372
rect 529934 21360 529940 21372
rect 529992 21360 529998 21412
rect 456702 20000 456708 20052
rect 456760 20040 456766 20052
rect 516134 20040 516140 20052
rect 456760 20012 516140 20040
rect 456760 20000 456766 20012
rect 516134 20000 516140 20012
rect 516192 20000 516198 20052
rect 75822 19932 75828 19984
rect 75880 19972 75886 19984
rect 136634 19972 136640 19984
rect 75880 19944 136640 19972
rect 75880 19932 75886 19944
rect 136634 19932 136640 19944
rect 136692 19932 136698 19984
rect 140682 19932 140688 19984
rect 140740 19972 140746 19984
rect 201586 19972 201592 19984
rect 140740 19944 201592 19972
rect 140740 19932 140746 19944
rect 201586 19932 201592 19944
rect 201644 19932 201650 19984
rect 208302 19932 208308 19984
rect 208360 19972 208366 19984
rect 269114 19972 269120 19984
rect 208360 19944 269120 19972
rect 208360 19932 208366 19944
rect 269114 19932 269120 19944
rect 269172 19932 269178 19984
rect 273162 19932 273168 19984
rect 273220 19972 273226 19984
rect 332594 19972 332600 19984
rect 273220 19944 332600 19972
rect 273220 19932 273226 19944
rect 332594 19932 332600 19944
rect 332652 19932 332658 19984
rect 333882 19932 333888 19984
rect 333940 19972 333946 19984
rect 393314 19972 393320 19984
rect 333940 19944 393320 19972
rect 333940 19932 333946 19944
rect 393314 19932 393320 19944
rect 393372 19932 393378 19984
rect 405642 19932 405648 19984
rect 405700 19972 405706 19984
rect 465074 19972 465080 19984
rect 405700 19944 465080 19972
rect 405700 19932 405706 19944
rect 465074 19932 465080 19944
rect 465132 19932 465138 19984
rect 506382 19932 506388 19984
rect 506440 19972 506446 19984
rect 565814 19972 565820 19984
rect 506440 19944 565820 19972
rect 506440 19932 506446 19944
rect 565814 19932 565820 19944
rect 565872 19932 565878 19984
rect 412634 19360 412640 19372
rect 412595 19332 412640 19360
rect 412634 19320 412640 19332
rect 412692 19320 412698 19372
rect 372614 19292 372620 19304
rect 372575 19264 372620 19292
rect 372614 19252 372620 19264
rect 372672 19252 372678 19304
rect 390370 19252 390376 19304
rect 390428 19292 390434 19304
rect 390554 19292 390560 19304
rect 390428 19264 390560 19292
rect 390428 19252 390434 19264
rect 390554 19252 390560 19264
rect 390612 19252 390618 19304
rect 434806 19292 434812 19304
rect 434767 19264 434812 19292
rect 434806 19252 434812 19264
rect 434864 19252 434870 19304
rect 467098 18640 467104 18692
rect 467156 18680 467162 18692
rect 520366 18680 520372 18692
rect 467156 18652 520372 18680
rect 467156 18640 467162 18652
rect 520366 18640 520372 18652
rect 520424 18640 520430 18692
rect 73062 18572 73068 18624
rect 73120 18612 73126 18624
rect 132586 18612 132592 18624
rect 73120 18584 132592 18612
rect 73120 18572 73126 18584
rect 132586 18572 132592 18584
rect 132644 18572 132650 18624
rect 136450 18572 136456 18624
rect 136508 18612 136514 18624
rect 197354 18612 197360 18624
rect 136508 18584 197360 18612
rect 136508 18572 136514 18584
rect 197354 18572 197360 18584
rect 197412 18572 197418 18624
rect 201402 18572 201408 18624
rect 201460 18612 201466 18624
rect 262306 18612 262312 18624
rect 201460 18584 262312 18612
rect 201460 18572 201466 18584
rect 262306 18572 262312 18584
rect 262364 18572 262370 18624
rect 266262 18572 266268 18624
rect 266320 18612 266326 18624
rect 325694 18612 325700 18624
rect 266320 18584 325700 18612
rect 266320 18572 266326 18584
rect 325694 18572 325700 18584
rect 325752 18572 325758 18624
rect 326982 18572 326988 18624
rect 327040 18612 327046 18624
rect 386414 18612 386420 18624
rect 327040 18584 386420 18612
rect 327040 18572 327046 18584
rect 386414 18572 386420 18584
rect 386472 18572 386478 18624
rect 408402 18572 408408 18624
rect 408460 18612 408466 18624
rect 467834 18612 467840 18624
rect 408460 18584 467840 18612
rect 408460 18572 408466 18584
rect 467834 18572 467840 18584
rect 467892 18572 467898 18624
rect 510522 18572 510528 18624
rect 510580 18612 510586 18624
rect 569954 18612 569960 18624
rect 510580 18584 569960 18612
rect 510580 18572 510586 18584
rect 569954 18572 569960 18584
rect 570012 18572 570018 18624
rect 523770 17892 523776 17944
rect 523828 17932 523834 17944
rect 580074 17932 580080 17944
rect 523828 17904 580080 17932
rect 523828 17892 523834 17904
rect 580074 17892 580080 17904
rect 580132 17892 580138 17944
rect 70302 17280 70308 17332
rect 70360 17320 70366 17332
rect 131114 17320 131120 17332
rect 70360 17292 131120 17320
rect 70360 17280 70366 17292
rect 131114 17280 131120 17292
rect 131172 17280 131178 17332
rect 401502 17280 401508 17332
rect 401560 17320 401566 17332
rect 460934 17320 460940 17332
rect 401560 17292 460940 17320
rect 401560 17280 401566 17292
rect 460934 17280 460940 17292
rect 460992 17280 460998 17332
rect 129642 17212 129648 17264
rect 129700 17252 129706 17264
rect 190454 17252 190460 17264
rect 129700 17224 190460 17252
rect 129700 17212 129706 17224
rect 190454 17212 190460 17224
rect 190512 17212 190518 17264
rect 197170 17212 197176 17264
rect 197228 17252 197234 17264
rect 258074 17252 258080 17264
rect 197228 17224 258080 17252
rect 197228 17212 197234 17224
rect 258074 17212 258080 17224
rect 258132 17212 258138 17264
rect 262122 17212 262128 17264
rect 262180 17252 262186 17264
rect 321646 17252 321652 17264
rect 262180 17224 321652 17252
rect 262180 17212 262186 17224
rect 321646 17212 321652 17224
rect 321704 17212 321710 17264
rect 322842 17212 322848 17264
rect 322900 17252 322906 17264
rect 382366 17252 382372 17264
rect 322900 17224 382372 17252
rect 322900 17212 322906 17224
rect 382366 17212 382372 17224
rect 382424 17212 382430 17264
rect 452562 17212 452568 17264
rect 452620 17252 452626 17264
rect 512086 17252 512092 17264
rect 452620 17224 512092 17252
rect 452620 17212 452626 17224
rect 512086 17212 512092 17224
rect 512144 17212 512150 17264
rect 126790 15920 126796 15972
rect 126848 15960 126854 15972
rect 186314 15960 186320 15972
rect 126848 15932 186320 15960
rect 126848 15920 126854 15932
rect 186314 15920 186320 15932
rect 186372 15920 186378 15972
rect 315942 15920 315948 15972
rect 316000 15960 316006 15972
rect 375374 15960 375380 15972
rect 316000 15932 375380 15960
rect 316000 15920 316006 15932
rect 375374 15920 375380 15932
rect 375432 15920 375438 15972
rect 424962 15920 424968 15972
rect 425020 15960 425026 15972
rect 485774 15960 485780 15972
rect 425020 15932 485780 15960
rect 425020 15920 425026 15932
rect 485774 15920 485780 15932
rect 485832 15920 485838 15972
rect 66898 15852 66904 15904
rect 66956 15892 66962 15904
rect 126974 15892 126980 15904
rect 66956 15864 126980 15892
rect 66956 15852 66962 15864
rect 126974 15852 126980 15864
rect 127032 15852 127038 15904
rect 194502 15852 194508 15904
rect 194560 15892 194566 15904
rect 253934 15892 253940 15904
rect 194560 15864 253940 15892
rect 194560 15852 194566 15864
rect 253934 15852 253940 15864
rect 253992 15852 253998 15904
rect 257890 15852 257896 15904
rect 257948 15892 257954 15904
rect 318794 15892 318800 15904
rect 257948 15864 318800 15892
rect 257948 15852 257954 15864
rect 318794 15852 318800 15864
rect 318852 15852 318858 15904
rect 397362 15852 397368 15904
rect 397420 15892 397426 15904
rect 458174 15892 458180 15904
rect 397420 15864 458180 15892
rect 397420 15852 397426 15864
rect 458174 15852 458180 15864
rect 458232 15852 458238 15904
rect 469122 15852 469128 15904
rect 469180 15892 469186 15904
rect 528646 15892 528652 15904
rect 469180 15864 528652 15892
rect 469180 15852 469186 15864
rect 528646 15852 528652 15864
rect 528704 15852 528710 15904
rect 81342 14492 81348 14544
rect 81400 14532 81406 14544
rect 140866 14532 140872 14544
rect 81400 14504 140872 14532
rect 81400 14492 81406 14504
rect 140866 14492 140872 14504
rect 140924 14492 140930 14544
rect 309042 14492 309048 14544
rect 309100 14532 309106 14544
rect 368474 14532 368480 14544
rect 309100 14504 368480 14532
rect 309100 14492 309106 14504
rect 368474 14492 368480 14504
rect 368532 14492 368538 14544
rect 395982 14492 395988 14544
rect 396040 14532 396046 14544
rect 455414 14532 455420 14544
rect 396040 14504 455420 14532
rect 396040 14492 396046 14504
rect 455414 14492 455420 14504
rect 455472 14492 455478 14544
rect 122742 14424 122748 14476
rect 122800 14464 122806 14476
rect 183646 14464 183652 14476
rect 122800 14436 183652 14464
rect 122800 14424 122806 14436
rect 183646 14424 183652 14436
rect 183704 14424 183710 14476
rect 187602 14424 187608 14476
rect 187660 14464 187666 14476
rect 247034 14464 247040 14476
rect 187660 14436 247040 14464
rect 187660 14424 187666 14436
rect 247034 14424 247040 14436
rect 247092 14424 247098 14476
rect 251082 14424 251088 14476
rect 251140 14464 251146 14476
rect 311894 14464 311900 14476
rect 251140 14436 311900 14464
rect 251140 14424 251146 14436
rect 311894 14424 311900 14436
rect 311952 14424 311958 14476
rect 344922 14424 344928 14476
rect 344980 14464 344986 14476
rect 405734 14464 405740 14476
rect 344980 14436 405740 14464
rect 344980 14424 344986 14436
rect 405734 14424 405740 14436
rect 405792 14424 405798 14476
rect 448422 14424 448428 14476
rect 448480 14464 448486 14476
rect 507854 14464 507860 14476
rect 448480 14436 507860 14464
rect 448480 14424 448486 14436
rect 507854 14424 507860 14436
rect 507912 14424 507918 14476
rect 509142 14424 509148 14476
rect 509200 14464 509206 14476
rect 568574 14464 568580 14476
rect 509200 14436 568580 14464
rect 509200 14424 509206 14436
rect 568574 14424 568580 14436
rect 568632 14424 568638 14476
rect 84102 13132 84108 13184
rect 84160 13172 84166 13184
rect 144914 13172 144920 13184
rect 84160 13144 144920 13172
rect 84160 13132 84166 13144
rect 144914 13132 144920 13144
rect 144972 13132 144978 13184
rect 248322 13132 248328 13184
rect 248380 13172 248386 13184
rect 307754 13172 307760 13184
rect 248380 13144 307760 13172
rect 248380 13132 248386 13144
rect 307754 13132 307760 13144
rect 307812 13132 307818 13184
rect 367738 13132 367744 13184
rect 367796 13172 367802 13184
rect 394694 13172 394700 13184
rect 367796 13144 394700 13172
rect 367796 13132 367802 13144
rect 394694 13132 394700 13144
rect 394752 13132 394758 13184
rect 444282 13132 444288 13184
rect 444340 13172 444346 13184
rect 503714 13172 503720 13184
rect 444340 13144 503720 13172
rect 444340 13132 444346 13144
rect 503714 13132 503720 13144
rect 503772 13132 503778 13184
rect 118510 13064 118516 13116
rect 118568 13104 118574 13116
rect 179414 13104 179420 13116
rect 118568 13076 179420 13104
rect 118568 13064 118574 13076
rect 179414 13064 179420 13076
rect 179472 13064 179478 13116
rect 183462 13064 183468 13116
rect 183520 13104 183526 13116
rect 244366 13104 244372 13116
rect 183520 13076 244372 13104
rect 183520 13064 183526 13076
rect 244366 13064 244372 13076
rect 244424 13064 244430 13116
rect 304902 13064 304908 13116
rect 304960 13104 304966 13116
rect 365806 13104 365812 13116
rect 304960 13076 365812 13104
rect 304960 13064 304966 13076
rect 365806 13064 365812 13076
rect 365864 13064 365870 13116
rect 389082 13064 389088 13116
rect 389140 13104 389146 13116
rect 448514 13104 448520 13116
rect 389140 13076 448520 13104
rect 389140 13064 389146 13076
rect 448514 13064 448520 13076
rect 448572 13064 448578 13116
rect 505002 13064 505008 13116
rect 505060 13104 505066 13116
rect 564434 13104 564440 13116
rect 505060 13076 564440 13104
rect 505060 13064 505066 13076
rect 564434 13064 564440 13076
rect 564492 13064 564498 13116
rect 383286 12384 383292 12436
rect 383344 12424 383350 12436
rect 383470 12424 383476 12436
rect 383344 12396 383476 12424
rect 383344 12384 383350 12396
rect 383470 12384 383476 12396
rect 383528 12384 383534 12436
rect 401594 12384 401600 12436
rect 401652 12424 401658 12436
rect 402514 12424 402520 12436
rect 401652 12396 402520 12424
rect 401652 12384 401658 12396
rect 402514 12384 402520 12396
rect 402572 12384 402578 12436
rect 404354 12384 404360 12436
rect 404412 12424 404418 12436
rect 404906 12424 404912 12436
rect 404412 12396 404912 12424
rect 404412 12384 404418 12396
rect 404906 12384 404912 12396
rect 404964 12384 404970 12436
rect 372617 12291 372675 12297
rect 372617 12257 372629 12291
rect 372663 12288 372675 12291
rect 372798 12288 372804 12300
rect 372663 12260 372804 12288
rect 372663 12257 372675 12260
rect 372617 12251 372675 12257
rect 372798 12248 372804 12260
rect 372856 12248 372862 12300
rect 331122 11772 331128 11824
rect 331180 11812 331186 11824
rect 391842 11812 391848 11824
rect 331180 11784 391848 11812
rect 331180 11772 331186 11784
rect 391842 11772 391848 11784
rect 391900 11772 391906 11824
rect 441522 11772 441528 11824
rect 441580 11812 441586 11824
rect 500954 11812 500960 11824
rect 441580 11784 500960 11812
rect 441580 11772 441586 11784
rect 500954 11772 500960 11784
rect 501012 11772 501018 11824
rect 115842 11704 115848 11756
rect 115900 11744 115906 11756
rect 175366 11744 175372 11756
rect 115900 11716 175372 11744
rect 115900 11704 115906 11716
rect 175366 11704 175372 11716
rect 175424 11704 175430 11756
rect 179230 11704 179236 11756
rect 179288 11744 179294 11756
rect 240134 11744 240140 11756
rect 179288 11716 240140 11744
rect 179288 11704 179294 11716
rect 240134 11704 240140 11716
rect 240192 11704 240198 11756
rect 241422 11704 241428 11756
rect 241480 11744 241486 11756
rect 300854 11744 300860 11756
rect 241480 11716 300860 11744
rect 241480 11704 241486 11716
rect 300854 11704 300860 11716
rect 300912 11704 300918 11756
rect 302142 11704 302148 11756
rect 302200 11744 302206 11756
rect 361574 11744 361580 11756
rect 302200 11716 361580 11744
rect 302200 11704 302206 11716
rect 361574 11704 361580 11716
rect 361632 11704 361638 11756
rect 380710 11704 380716 11756
rect 380768 11744 380774 11756
rect 441614 11744 441620 11756
rect 380768 11716 441620 11744
rect 380768 11704 380774 11716
rect 441614 11704 441620 11716
rect 441672 11704 441678 11756
rect 499482 11704 499488 11756
rect 499540 11744 499546 11756
rect 558914 11744 558920 11756
rect 499540 11716 558920 11744
rect 499540 11704 499546 11716
rect 558914 11704 558920 11716
rect 558972 11704 558978 11756
rect 311158 10412 311164 10464
rect 311216 10452 311222 10464
rect 370406 10452 370412 10464
rect 311216 10424 370412 10452
rect 311216 10412 311222 10424
rect 370406 10412 370412 10424
rect 370464 10412 370470 10464
rect 176562 10344 176568 10396
rect 176620 10384 176626 10396
rect 236086 10384 236092 10396
rect 176620 10356 236092 10384
rect 176620 10344 176626 10356
rect 236086 10344 236092 10356
rect 236144 10344 236150 10396
rect 298002 10344 298008 10396
rect 298060 10384 298066 10396
rect 357434 10384 357440 10396
rect 298060 10356 357440 10384
rect 298060 10344 298066 10356
rect 357434 10344 357440 10356
rect 357492 10344 357498 10396
rect 416682 10344 416688 10396
rect 416740 10384 416746 10396
rect 477586 10384 477592 10396
rect 416740 10356 477592 10384
rect 416740 10344 416746 10356
rect 477586 10344 477592 10356
rect 477644 10344 477650 10396
rect 111702 10276 111708 10328
rect 111760 10316 111766 10328
rect 172514 10316 172520 10328
rect 111760 10288 172520 10316
rect 111760 10276 111766 10288
rect 172514 10276 172520 10288
rect 172572 10276 172578 10328
rect 233142 10276 233148 10328
rect 233200 10316 233206 10328
rect 293954 10316 293960 10328
rect 233200 10288 293960 10316
rect 233200 10276 233206 10288
rect 293954 10276 293960 10288
rect 294012 10276 294018 10328
rect 355962 10276 355968 10328
rect 356020 10316 356026 10328
rect 416866 10316 416872 10328
rect 356020 10288 416872 10316
rect 356020 10276 356026 10288
rect 416866 10276 416872 10288
rect 416924 10276 416930 10328
rect 437382 10276 437388 10328
rect 437440 10316 437446 10328
rect 496814 10316 496820 10328
rect 437440 10288 496820 10316
rect 437440 10276 437446 10288
rect 496814 10276 496820 10288
rect 496872 10276 496878 10328
rect 498102 10276 498108 10328
rect 498160 10316 498166 10328
rect 557534 10316 557540 10328
rect 498160 10288 557540 10316
rect 498160 10276 498166 10288
rect 557534 10276 557540 10288
rect 557592 10276 557598 10328
rect 434806 9772 434812 9784
rect 434767 9744 434812 9772
rect 434806 9732 434812 9744
rect 434864 9732 434870 9784
rect 390646 9596 390652 9648
rect 390704 9596 390710 9648
rect 411254 9596 411260 9648
rect 411312 9636 411318 9648
rect 412085 9639 412143 9645
rect 412085 9636 412097 9639
rect 411312 9608 412097 9636
rect 411312 9596 411318 9608
rect 412085 9605 412097 9608
rect 412131 9605 412143 9639
rect 412085 9599 412143 9605
rect 415394 9596 415400 9648
rect 415452 9636 415458 9648
rect 415673 9639 415731 9645
rect 415673 9636 415685 9639
rect 415452 9608 415685 9636
rect 415452 9596 415458 9608
rect 415673 9605 415685 9608
rect 415719 9605 415731 9639
rect 415673 9599 415731 9605
rect 434806 9596 434812 9648
rect 434864 9636 434870 9648
rect 435821 9639 435879 9645
rect 435821 9636 435833 9639
rect 434864 9608 435833 9636
rect 434864 9596 434870 9608
rect 435821 9605 435833 9608
rect 435867 9605 435879 9639
rect 435821 9599 435879 9605
rect 390664 9512 390692 9596
rect 390646 9460 390652 9512
rect 390704 9460 390710 9512
rect 230382 8984 230388 9036
rect 230440 9024 230446 9036
rect 290734 9024 290740 9036
rect 230440 8996 290740 9024
rect 230440 8984 230446 8996
rect 290734 8984 290740 8996
rect 290792 8984 290798 9036
rect 291102 8984 291108 9036
rect 291160 9024 291166 9036
rect 351362 9024 351368 9036
rect 291160 8996 351368 9024
rect 291160 8984 291166 8996
rect 351362 8984 351368 8996
rect 351420 8984 351426 9036
rect 108942 8916 108948 8968
rect 109000 8956 109006 8968
rect 169386 8956 169392 8968
rect 109000 8928 169392 8956
rect 109000 8916 109006 8928
rect 169386 8916 169392 8928
rect 169444 8916 169450 8968
rect 172422 8916 172428 8968
rect 172480 8956 172486 8968
rect 233694 8956 233700 8968
rect 172480 8928 233700 8956
rect 172480 8916 172486 8928
rect 233694 8916 233700 8928
rect 233752 8916 233758 8968
rect 347682 8916 347688 8968
rect 347740 8956 347746 8968
rect 408586 8956 408592 8968
rect 347740 8928 408592 8956
rect 347740 8916 347746 8928
rect 408586 8916 408592 8928
rect 408644 8916 408650 8968
rect 430482 8916 430488 8968
rect 430540 8956 430546 8968
rect 490558 8956 490564 8968
rect 430540 8928 490564 8956
rect 430540 8916 430546 8928
rect 490558 8916 490564 8928
rect 490616 8916 490622 8968
rect 491202 8916 491208 8968
rect 491260 8956 491266 8968
rect 551186 8956 551192 8968
rect 491260 8928 551192 8956
rect 491260 8916 491266 8928
rect 551186 8916 551192 8928
rect 551244 8916 551250 8968
rect 137922 7624 137928 7676
rect 137980 7664 137986 7676
rect 199194 7664 199200 7676
rect 137980 7636 199200 7664
rect 137980 7624 137986 7636
rect 199194 7624 199200 7636
rect 199252 7624 199258 7676
rect 223482 7624 223488 7676
rect 223540 7664 223546 7676
rect 283650 7664 283656 7676
rect 223540 7636 283656 7664
rect 223540 7624 223546 7636
rect 283650 7624 283656 7636
rect 283708 7624 283714 7676
rect 340782 7624 340788 7676
rect 340840 7664 340846 7676
rect 401318 7664 401324 7676
rect 340840 7636 401324 7664
rect 340840 7624 340846 7636
rect 401318 7624 401324 7636
rect 401376 7624 401382 7676
rect 433334 7624 433340 7676
rect 433392 7664 433398 7676
rect 434622 7664 434628 7676
rect 433392 7636 434628 7664
rect 433392 7624 433398 7636
rect 434622 7624 434628 7636
rect 434680 7624 434686 7676
rect 481542 7624 481548 7676
rect 481600 7664 481606 7676
rect 541710 7664 541716 7676
rect 481600 7636 541716 7664
rect 481600 7624 481606 7636
rect 541710 7624 541716 7636
rect 541768 7624 541774 7676
rect 104802 7556 104808 7608
rect 104860 7596 104866 7608
rect 165890 7596 165896 7608
rect 104860 7568 165896 7596
rect 104860 7556 104866 7568
rect 165890 7556 165896 7568
rect 165948 7556 165954 7608
rect 169662 7556 169668 7608
rect 169720 7596 169726 7608
rect 230106 7596 230112 7608
rect 169720 7568 230112 7596
rect 169720 7556 169726 7568
rect 230106 7556 230112 7568
rect 230164 7556 230170 7608
rect 284202 7556 284208 7608
rect 284260 7596 284266 7608
rect 344278 7596 344284 7608
rect 284260 7568 344284 7596
rect 284260 7556 284266 7568
rect 344278 7556 344284 7568
rect 344336 7556 344342 7608
rect 382366 7556 382372 7608
rect 382424 7596 382430 7608
rect 383562 7596 383568 7608
rect 382424 7568 383568 7596
rect 382424 7556 382430 7568
rect 383562 7556 383568 7568
rect 383620 7556 383626 7608
rect 408494 7556 408500 7608
rect 408552 7596 408558 7608
rect 409690 7596 409696 7608
rect 408552 7568 409696 7596
rect 408552 7556 408558 7568
rect 409690 7556 409696 7568
rect 409748 7556 409754 7608
rect 426342 7556 426348 7608
rect 426400 7596 426406 7608
rect 486970 7596 486976 7608
rect 426400 7568 486976 7596
rect 426400 7556 426406 7568
rect 486970 7556 486976 7568
rect 487028 7556 487034 7608
rect 162762 6264 162768 6316
rect 162820 6304 162826 6316
rect 222930 6304 222936 6316
rect 162820 6276 222936 6304
rect 162820 6264 162826 6276
rect 222930 6264 222936 6276
rect 222988 6264 222994 6316
rect 219342 6196 219348 6248
rect 219400 6236 219406 6248
rect 279970 6236 279976 6248
rect 219400 6208 279976 6236
rect 219400 6196 219406 6208
rect 279970 6196 279976 6208
rect 280028 6196 280034 6248
rect 282822 6196 282828 6248
rect 282880 6236 282886 6248
rect 343082 6236 343088 6248
rect 282880 6208 343088 6236
rect 282880 6196 282886 6208
rect 343082 6196 343088 6208
rect 343140 6196 343146 6248
rect 423582 6196 423588 6248
rect 423640 6236 423646 6248
rect 483474 6236 483480 6248
rect 423640 6208 483480 6236
rect 423640 6196 423646 6208
rect 483474 6196 483480 6208
rect 483532 6196 483538 6248
rect 100570 6128 100576 6180
rect 100628 6168 100634 6180
rect 162302 6168 162308 6180
rect 100628 6140 162308 6168
rect 100628 6128 100634 6140
rect 162302 6128 162308 6140
rect 162360 6128 162366 6180
rect 209682 6128 209688 6180
rect 209740 6168 209746 6180
rect 270586 6168 270592 6180
rect 209740 6140 270592 6168
rect 209740 6128 209746 6140
rect 270586 6128 270592 6140
rect 270644 6128 270650 6180
rect 280062 6128 280068 6180
rect 280120 6168 280126 6180
rect 340690 6168 340696 6180
rect 280120 6140 340696 6168
rect 280120 6128 280126 6140
rect 340690 6128 340696 6140
rect 340748 6128 340754 6180
rect 345658 6128 345664 6180
rect 345716 6168 345722 6180
rect 379974 6168 379980 6180
rect 345716 6140 379980 6168
rect 345716 6128 345722 6140
rect 379974 6128 379980 6140
rect 380032 6128 380038 6180
rect 398742 6128 398748 6180
rect 398800 6168 398806 6180
rect 459646 6168 459652 6180
rect 398800 6140 459652 6168
rect 398800 6128 398806 6140
rect 459646 6128 459652 6140
rect 459704 6128 459710 6180
rect 516042 6128 516048 6180
rect 516100 6168 516106 6180
rect 576210 6168 576216 6180
rect 516100 6140 576216 6168
rect 516100 6128 516106 6140
rect 576210 6128 576216 6140
rect 576268 6128 576274 6180
rect 380802 5448 380808 5500
rect 380860 5488 380866 5500
rect 440602 5488 440608 5500
rect 380860 5460 440608 5488
rect 380860 5448 380866 5460
rect 440602 5448 440608 5460
rect 440660 5448 440666 5500
rect 369762 5380 369768 5432
rect 369820 5420 369826 5432
rect 429930 5420 429936 5432
rect 369820 5392 429936 5420
rect 369820 5380 369826 5392
rect 429930 5380 429936 5392
rect 429988 5380 429994 5432
rect 455322 5380 455328 5432
rect 455380 5420 455386 5432
rect 515582 5420 515588 5432
rect 455380 5392 515588 5420
rect 455380 5380 455386 5392
rect 515582 5380 515588 5392
rect 515640 5380 515646 5432
rect 365622 5312 365628 5364
rect 365680 5352 365686 5364
rect 426342 5352 426348 5364
rect 365680 5324 426348 5352
rect 365680 5312 365686 5324
rect 426342 5312 426348 5324
rect 426400 5312 426406 5364
rect 459462 5312 459468 5364
rect 459520 5352 459526 5364
rect 519078 5352 519084 5364
rect 459520 5324 519084 5352
rect 459520 5312 459526 5324
rect 519078 5312 519084 5324
rect 519136 5312 519142 5364
rect 387702 5244 387708 5296
rect 387760 5284 387766 5296
rect 447778 5284 447784 5296
rect 387760 5256 447784 5284
rect 387760 5244 387766 5256
rect 447778 5244 447784 5256
rect 447836 5244 447842 5296
rect 462222 5244 462228 5296
rect 462280 5284 462286 5296
rect 522666 5284 522672 5296
rect 462280 5256 522672 5284
rect 462280 5244 462286 5256
rect 522666 5244 522672 5256
rect 522724 5244 522730 5296
rect 376662 5176 376668 5228
rect 376720 5216 376726 5228
rect 437014 5216 437020 5228
rect 376720 5188 437020 5216
rect 376720 5176 376726 5188
rect 437014 5176 437020 5188
rect 437072 5176 437078 5228
rect 466362 5176 466368 5228
rect 466420 5216 466426 5228
rect 526254 5216 526260 5228
rect 466420 5188 526260 5216
rect 466420 5176 466426 5188
rect 526254 5176 526260 5188
rect 526312 5176 526318 5228
rect 358722 5108 358728 5160
rect 358780 5148 358786 5160
rect 419166 5148 419172 5160
rect 358780 5120 419172 5148
rect 358780 5108 358786 5120
rect 419166 5108 419172 5120
rect 419224 5108 419230 5160
rect 473262 5108 473268 5160
rect 473320 5148 473326 5160
rect 533430 5148 533436 5160
rect 473320 5120 533436 5148
rect 473320 5108 473326 5120
rect 533430 5108 533436 5120
rect 533488 5108 533494 5160
rect 394602 5040 394608 5092
rect 394660 5080 394666 5092
rect 454862 5080 454868 5092
rect 394660 5052 454868 5080
rect 394660 5040 394666 5052
rect 454862 5040 454868 5052
rect 454920 5040 454926 5092
rect 480162 5040 480168 5092
rect 480220 5080 480226 5092
rect 540514 5080 540520 5092
rect 480220 5052 540520 5080
rect 480220 5040 480226 5052
rect 540514 5040 540520 5052
rect 540572 5040 540578 5092
rect 362862 4972 362868 5024
rect 362920 5012 362926 5024
rect 422754 5012 422760 5024
rect 362920 4984 422760 5012
rect 362920 4972 362926 4984
rect 422754 4972 422760 4984
rect 422812 4972 422818 5024
rect 484302 4972 484308 5024
rect 484360 5012 484366 5024
rect 544102 5012 544108 5024
rect 484360 4984 544108 5012
rect 484360 4972 484366 4984
rect 544102 4972 544108 4984
rect 544160 4972 544166 5024
rect 133782 4904 133788 4956
rect 133840 4944 133846 4956
rect 194410 4944 194416 4956
rect 133840 4916 194416 4944
rect 133840 4904 133846 4916
rect 194410 4904 194416 4916
rect 194468 4904 194474 4956
rect 255222 4904 255228 4956
rect 255280 4944 255286 4956
rect 315758 4944 315764 4956
rect 255280 4916 315764 4944
rect 255280 4904 255286 4916
rect 315758 4904 315764 4916
rect 315816 4904 315822 4956
rect 383286 4904 383292 4956
rect 383344 4944 383350 4956
rect 444190 4944 444196 4956
rect 383344 4916 444196 4944
rect 383344 4904 383350 4916
rect 444190 4904 444196 4916
rect 444248 4904 444254 4956
rect 463602 4904 463608 4956
rect 463660 4944 463666 4956
rect 523862 4944 523868 4956
rect 463660 4916 523868 4944
rect 463660 4904 463666 4916
rect 523862 4904 523868 4916
rect 523920 4904 523926 4956
rect 66162 4836 66168 4888
rect 66220 4876 66226 4888
rect 126606 4876 126612 4888
rect 66220 4848 126612 4876
rect 66220 4836 66226 4848
rect 126606 4836 126612 4848
rect 126664 4836 126670 4888
rect 190362 4836 190368 4888
rect 190420 4876 190426 4888
rect 251450 4876 251456 4888
rect 190420 4848 251456 4876
rect 190420 4836 190426 4848
rect 251450 4836 251456 4848
rect 251508 4836 251514 4888
rect 303522 4836 303528 4888
rect 303580 4876 303586 4888
rect 364518 4876 364524 4888
rect 303580 4848 364524 4876
rect 303580 4836 303586 4848
rect 364518 4836 364524 4848
rect 364576 4836 364582 4888
rect 390462 4836 390468 4888
rect 390520 4876 390526 4888
rect 396077 4879 396135 4885
rect 396077 4876 396089 4879
rect 390520 4848 396089 4876
rect 390520 4836 390526 4848
rect 396077 4845 396089 4848
rect 396123 4845 396135 4879
rect 396077 4839 396135 4845
rect 405737 4879 405795 4885
rect 405737 4845 405749 4879
rect 405783 4845 405795 4879
rect 405737 4839 405795 4845
rect 413281 4879 413339 4885
rect 413281 4845 413293 4879
rect 413327 4876 413339 4879
rect 422941 4879 422999 4885
rect 422941 4876 422953 4879
rect 413327 4848 422953 4876
rect 413327 4845 413339 4848
rect 413281 4839 413339 4845
rect 422941 4845 422953 4848
rect 422987 4845 422999 4879
rect 422941 4839 422999 4845
rect 427817 4879 427875 4885
rect 427817 4845 427829 4879
rect 427863 4876 427875 4879
rect 427863 4848 446444 4876
rect 427863 4845 427875 4848
rect 427817 4839 427875 4845
rect 68922 4768 68928 4820
rect 68980 4808 68986 4820
rect 130194 4808 130200 4820
rect 68980 4780 130200 4808
rect 68980 4768 68986 4780
rect 130194 4768 130200 4780
rect 130252 4768 130258 4820
rect 173802 4768 173808 4820
rect 173860 4808 173866 4820
rect 234798 4808 234804 4820
rect 173860 4780 234804 4808
rect 173860 4768 173866 4780
rect 234798 4768 234804 4780
rect 234856 4768 234862 4820
rect 252462 4768 252468 4820
rect 252520 4808 252526 4820
rect 313366 4808 313372 4820
rect 252520 4780 313372 4808
rect 252520 4768 252526 4780
rect 313366 4768 313372 4780
rect 313424 4768 313430 4820
rect 372522 4768 372528 4820
rect 372580 4808 372586 4820
rect 395985 4811 396043 4817
rect 372580 4780 379560 4808
rect 372580 4768 372586 4780
rect 379532 4740 379560 4780
rect 395985 4777 395997 4811
rect 396031 4808 396043 4811
rect 405752 4808 405780 4839
rect 425054 4808 425060 4820
rect 396031 4780 405780 4808
rect 418172 4780 425060 4808
rect 396031 4777 396043 4780
rect 395985 4771 396043 4777
rect 396077 4743 396135 4749
rect 379532 4712 390324 4740
rect 390296 4672 390324 4712
rect 396077 4709 396089 4743
rect 396123 4740 396135 4743
rect 405737 4743 405795 4749
rect 396123 4712 396580 4740
rect 396123 4709 396135 4712
rect 396077 4703 396135 4709
rect 395985 4675 396043 4681
rect 395985 4672 395997 4675
rect 390296 4644 395997 4672
rect 395985 4641 395997 4644
rect 396031 4641 396043 4675
rect 396552 4672 396580 4712
rect 405737 4709 405749 4743
rect 405783 4740 405795 4743
rect 405783 4712 418016 4740
rect 405783 4709 405795 4712
rect 405737 4703 405795 4709
rect 413281 4675 413339 4681
rect 413281 4672 413293 4675
rect 396552 4644 413293 4672
rect 395985 4635 396043 4641
rect 413281 4641 413293 4644
rect 413327 4641 413339 4675
rect 417988 4672 418016 4712
rect 418172 4672 418200 4780
rect 425054 4768 425060 4780
rect 425112 4768 425118 4820
rect 446416 4740 446444 4848
rect 487062 4836 487068 4888
rect 487120 4876 487126 4888
rect 547690 4876 547696 4888
rect 487120 4848 547696 4876
rect 487120 4836 487126 4848
rect 547690 4836 547696 4848
rect 547748 4836 547754 4888
rect 476022 4768 476028 4820
rect 476080 4808 476086 4820
rect 536926 4808 536932 4820
rect 476080 4780 536932 4808
rect 476080 4768 476086 4780
rect 536926 4768 536932 4780
rect 536984 4768 536990 4820
rect 451366 4740 451372 4752
rect 446416 4712 451372 4740
rect 451366 4700 451372 4712
rect 451424 4700 451430 4752
rect 417988 4644 418200 4672
rect 422941 4675 422999 4681
rect 413281 4635 413339 4641
rect 422941 4641 422953 4675
rect 422987 4672 422999 4675
rect 427725 4675 427783 4681
rect 427725 4672 427737 4675
rect 422987 4644 427737 4672
rect 422987 4641 422999 4644
rect 422941 4635 422999 4641
rect 427725 4641 427737 4644
rect 427771 4641 427783 4675
rect 427725 4635 427783 4641
rect 528646 4156 528652 4208
rect 528704 4196 528710 4208
rect 529842 4196 529848 4208
rect 528704 4168 529848 4196
rect 528704 4156 528710 4168
rect 529842 4156 529848 4168
rect 529900 4156 529906 4208
rect 118602 4088 118608 4140
rect 118660 4128 118666 4140
rect 178954 4128 178960 4140
rect 118660 4100 178960 4128
rect 118660 4088 118666 4100
rect 178954 4088 178960 4100
rect 179012 4088 179018 4140
rect 179322 4088 179328 4140
rect 179380 4128 179386 4140
rect 239582 4128 239588 4140
rect 179380 4100 239588 4128
rect 179380 4088 179386 4100
rect 239582 4088 239588 4100
rect 239640 4088 239646 4140
rect 264882 4088 264888 4140
rect 264940 4128 264946 4140
rect 325234 4128 325240 4140
rect 264940 4100 325240 4128
rect 264940 4088 264946 4100
rect 325234 4088 325240 4100
rect 325292 4088 325298 4140
rect 379422 4088 379428 4140
rect 379480 4128 379486 4140
rect 439406 4128 439412 4140
rect 379480 4100 439412 4128
rect 379480 4088 379486 4100
rect 439406 4088 439412 4100
rect 439464 4088 439470 4140
rect 442902 4088 442908 4140
rect 442960 4128 442966 4140
rect 503622 4128 503628 4140
rect 442960 4100 503628 4128
rect 442960 4088 442966 4100
rect 503622 4088 503628 4100
rect 503680 4088 503686 4140
rect 514662 4088 514668 4140
rect 514720 4128 514726 4140
rect 575014 4128 575020 4140
rect 514720 4100 575020 4128
rect 514720 4088 514726 4100
rect 575014 4088 575020 4100
rect 575072 4088 575078 4140
rect 150342 4020 150348 4072
rect 150400 4060 150406 4072
rect 211062 4060 211068 4072
rect 150400 4032 211068 4060
rect 150400 4020 150406 4032
rect 211062 4020 211068 4032
rect 211120 4020 211126 4072
rect 240042 4020 240048 4072
rect 240100 4060 240106 4072
rect 300302 4060 300308 4072
rect 240100 4032 300308 4060
rect 240100 4020 240106 4032
rect 300302 4020 300308 4032
rect 300360 4020 300366 4072
rect 350442 4020 350448 4072
rect 350500 4060 350506 4072
rect 410886 4060 410892 4072
rect 350500 4032 410892 4060
rect 350500 4020 350506 4032
rect 410886 4020 410892 4032
rect 410944 4020 410950 4072
rect 411162 4020 411168 4072
rect 411220 4060 411226 4072
rect 471514 4060 471520 4072
rect 411220 4032 471520 4060
rect 411220 4020 411226 4032
rect 471514 4020 471520 4032
rect 471572 4020 471578 4072
rect 493962 4020 493968 4072
rect 494020 4060 494026 4072
rect 553578 4060 553584 4072
rect 494020 4032 553584 4060
rect 494020 4020 494026 4032
rect 553578 4020 553584 4032
rect 553636 4020 553642 4072
rect 143442 3952 143448 4004
rect 143500 3992 143506 4004
rect 203886 3992 203892 4004
rect 143500 3964 203892 3992
rect 143500 3952 143506 3964
rect 203886 3952 203892 3964
rect 203944 3952 203950 4004
rect 231762 3952 231768 4004
rect 231820 3992 231826 4004
rect 237285 3995 237343 4001
rect 237285 3992 237297 3995
rect 231820 3964 237297 3992
rect 231820 3952 231826 3964
rect 237285 3961 237297 3964
rect 237331 3961 237343 3995
rect 237285 3955 237343 3961
rect 246942 3952 246948 4004
rect 247000 3992 247006 4004
rect 307386 3992 307392 4004
rect 247000 3964 307392 3992
rect 247000 3952 247006 3964
rect 307386 3952 307392 3964
rect 307444 3952 307450 4004
rect 318702 3952 318708 4004
rect 318760 3992 318766 4004
rect 378778 3992 378784 4004
rect 318760 3964 378784 3992
rect 318760 3952 318766 3964
rect 378778 3952 378784 3964
rect 378836 3952 378842 4004
rect 386322 3952 386328 4004
rect 386380 3992 386386 4004
rect 446582 3992 446588 4004
rect 386380 3964 446588 3992
rect 386380 3952 386386 3964
rect 446582 3952 446588 3964
rect 446640 3952 446646 4004
rect 496722 3952 496728 4004
rect 496780 3992 496786 4004
rect 557166 3992 557172 4004
rect 496780 3964 557172 3992
rect 496780 3952 496786 3964
rect 557166 3952 557172 3964
rect 557224 3952 557230 4004
rect 88242 3884 88248 3936
rect 88300 3924 88306 3936
rect 149238 3924 149244 3936
rect 88300 3896 149244 3924
rect 88300 3884 88306 3896
rect 149238 3884 149244 3896
rect 149296 3884 149302 3936
rect 161382 3884 161388 3936
rect 161440 3924 161446 3936
rect 221734 3924 221740 3936
rect 161440 3896 221740 3924
rect 161440 3884 161446 3896
rect 221734 3884 221740 3896
rect 221792 3884 221798 3936
rect 229002 3884 229008 3936
rect 229060 3924 229066 3936
rect 289538 3924 289544 3936
rect 229060 3896 289544 3924
rect 229060 3884 229066 3896
rect 289538 3884 289544 3896
rect 289596 3884 289602 3936
rect 300762 3884 300768 3936
rect 300820 3924 300826 3936
rect 360930 3924 360936 3936
rect 300820 3896 360936 3924
rect 300820 3884 300826 3896
rect 360930 3884 360936 3896
rect 360988 3884 360994 3936
rect 393222 3884 393228 3936
rect 393280 3924 393286 3936
rect 453666 3924 453672 3936
rect 393280 3896 453672 3924
rect 393280 3884 393286 3896
rect 453666 3884 453672 3896
rect 453724 3884 453730 3936
rect 500862 3884 500868 3936
rect 500920 3924 500926 3936
rect 560754 3924 560760 3936
rect 500920 3896 560760 3924
rect 500920 3884 500926 3896
rect 560754 3884 560760 3896
rect 560812 3884 560818 3936
rect 128262 3816 128268 3868
rect 128320 3856 128326 3868
rect 189626 3856 189632 3868
rect 128320 3828 189632 3856
rect 128320 3816 128326 3828
rect 189626 3816 189632 3828
rect 189684 3816 189690 3868
rect 197262 3816 197268 3868
rect 197320 3856 197326 3868
rect 257430 3856 257436 3868
rect 197320 3828 257436 3856
rect 197320 3816 197326 3828
rect 257430 3816 257436 3828
rect 257488 3816 257494 3868
rect 257982 3816 257988 3868
rect 258040 3856 258046 3868
rect 318058 3856 318064 3868
rect 258040 3828 318064 3856
rect 258040 3816 258046 3828
rect 318058 3816 318064 3828
rect 318116 3816 318122 3868
rect 325602 3816 325608 3868
rect 325660 3856 325666 3868
rect 385862 3856 385868 3868
rect 325660 3828 385868 3856
rect 325660 3816 325666 3828
rect 385862 3816 385868 3828
rect 385920 3816 385926 3868
rect 400122 3816 400128 3868
rect 400180 3856 400186 3868
rect 460750 3856 460756 3868
rect 400180 3828 460756 3856
rect 400180 3816 400186 3828
rect 460750 3816 460756 3828
rect 460808 3816 460814 3868
rect 503438 3816 503444 3868
rect 503496 3856 503502 3868
rect 564342 3856 564348 3868
rect 503496 3828 564348 3856
rect 503496 3816 503502 3828
rect 564342 3816 564348 3828
rect 564400 3816 564406 3868
rect 114462 3748 114468 3800
rect 114520 3788 114526 3800
rect 175274 3788 175280 3800
rect 114520 3760 175280 3788
rect 114520 3748 114526 3760
rect 175274 3748 175280 3760
rect 175332 3748 175338 3800
rect 200022 3748 200028 3800
rect 200080 3788 200086 3800
rect 261018 3788 261024 3800
rect 200080 3760 261024 3788
rect 200080 3748 200086 3760
rect 261018 3748 261024 3760
rect 261076 3748 261082 3800
rect 262214 3748 262220 3800
rect 262272 3788 262278 3800
rect 263410 3788 263416 3800
rect 262272 3760 263416 3788
rect 262272 3748 262278 3760
rect 263410 3748 263416 3760
rect 263468 3748 263474 3800
rect 289722 3748 289728 3800
rect 289780 3788 289786 3800
rect 350258 3788 350264 3800
rect 289780 3760 350264 3788
rect 289780 3748 289786 3760
rect 350258 3748 350264 3760
rect 350316 3748 350322 3800
rect 354582 3748 354588 3800
rect 354640 3788 354646 3800
rect 414474 3788 414480 3800
rect 354640 3760 414480 3788
rect 354640 3748 354646 3760
rect 414474 3748 414480 3760
rect 414532 3748 414538 3800
rect 447042 3748 447048 3800
rect 447100 3788 447106 3800
rect 507210 3788 507216 3800
rect 447100 3760 507216 3788
rect 447100 3748 447106 3760
rect 507210 3748 507216 3760
rect 507268 3748 507274 3800
rect 513282 3748 513288 3800
rect 513340 3788 513346 3800
rect 573818 3788 573824 3800
rect 513340 3760 573824 3788
rect 513340 3748 513346 3760
rect 573818 3748 573824 3760
rect 573876 3748 573882 3800
rect 121362 3680 121368 3732
rect 121420 3720 121426 3732
rect 182542 3720 182548 3732
rect 121420 3692 182548 3720
rect 121420 3680 121426 3692
rect 182542 3680 182548 3692
rect 182600 3680 182606 3732
rect 201494 3680 201500 3732
rect 201552 3720 201558 3732
rect 202690 3720 202696 3732
rect 201552 3692 202696 3720
rect 201552 3680 201558 3692
rect 202690 3680 202696 3692
rect 202748 3680 202754 3732
rect 206922 3680 206928 3732
rect 206980 3720 206986 3732
rect 268102 3720 268108 3732
rect 206980 3692 268108 3720
rect 206980 3680 206986 3692
rect 268102 3680 268108 3692
rect 268160 3680 268166 3732
rect 296622 3680 296628 3732
rect 296680 3720 296686 3732
rect 357342 3720 357348 3732
rect 296680 3692 357348 3720
rect 296680 3680 296686 3692
rect 357342 3680 357348 3692
rect 357400 3680 357406 3732
rect 361482 3680 361488 3732
rect 361540 3720 361546 3732
rect 421558 3720 421564 3732
rect 361540 3692 421564 3720
rect 361540 3680 361546 3692
rect 421558 3680 421564 3692
rect 421616 3680 421622 3732
rect 422202 3680 422208 3732
rect 422260 3720 422266 3732
rect 482278 3720 482284 3732
rect 422260 3692 482284 3720
rect 422260 3680 422266 3692
rect 482278 3680 482284 3692
rect 482336 3680 482342 3732
rect 511902 3680 511908 3732
rect 511960 3720 511966 3732
rect 571334 3720 571340 3732
rect 511960 3692 571340 3720
rect 511960 3680 511966 3692
rect 571334 3680 571340 3692
rect 571392 3680 571398 3732
rect 71682 3612 71688 3664
rect 71740 3652 71746 3664
rect 132494 3652 132500 3664
rect 71740 3624 132500 3652
rect 71740 3612 71746 3624
rect 132494 3612 132500 3624
rect 132552 3612 132558 3664
rect 153102 3612 153108 3664
rect 153160 3652 153166 3664
rect 214650 3652 214656 3664
rect 153160 3624 214656 3652
rect 153160 3612 153166 3624
rect 214650 3612 214656 3624
rect 214708 3612 214714 3664
rect 235902 3612 235908 3664
rect 235960 3652 235966 3664
rect 296714 3652 296720 3664
rect 235960 3624 296720 3652
rect 235960 3612 235966 3624
rect 296714 3612 296720 3624
rect 296772 3612 296778 3664
rect 321646 3612 321652 3664
rect 321704 3652 321710 3664
rect 322842 3652 322848 3664
rect 321704 3624 322848 3652
rect 321704 3612 321710 3624
rect 322842 3612 322848 3624
rect 322900 3612 322906 3664
rect 328362 3612 328368 3664
rect 328420 3652 328426 3664
rect 389450 3652 389456 3664
rect 328420 3624 389456 3652
rect 328420 3612 328426 3624
rect 389450 3612 389456 3624
rect 389508 3612 389514 3664
rect 418062 3612 418068 3664
rect 418120 3652 418126 3664
rect 478690 3652 478696 3664
rect 418120 3624 478696 3652
rect 418120 3612 418126 3624
rect 478690 3612 478696 3624
rect 478748 3612 478754 3664
rect 507762 3612 507768 3664
rect 507820 3652 507826 3664
rect 567838 3652 567844 3664
rect 507820 3624 567844 3652
rect 507820 3612 507826 3624
rect 567838 3612 567844 3624
rect 567896 3612 567902 3664
rect 78582 3544 78588 3596
rect 78640 3584 78646 3596
rect 139670 3584 139676 3596
rect 78640 3556 139676 3584
rect 78640 3544 78646 3556
rect 139670 3544 139676 3556
rect 139728 3544 139734 3596
rect 140866 3544 140872 3596
rect 140924 3584 140930 3596
rect 142062 3584 142068 3596
rect 140924 3556 142068 3584
rect 140924 3544 140930 3556
rect 142062 3544 142068 3556
rect 142120 3544 142126 3596
rect 150526 3544 150532 3596
rect 150584 3584 150590 3596
rect 151538 3584 151544 3596
rect 150584 3556 151544 3584
rect 150584 3544 150590 3556
rect 151538 3544 151544 3556
rect 151596 3544 151602 3596
rect 157242 3544 157248 3596
rect 157300 3584 157306 3596
rect 218054 3584 218060 3596
rect 157300 3556 218060 3584
rect 157300 3544 157306 3556
rect 218054 3544 218060 3556
rect 218112 3544 218118 3596
rect 218146 3544 218152 3596
rect 218204 3584 218210 3596
rect 219342 3584 219348 3596
rect 218204 3556 219348 3584
rect 218204 3544 218210 3556
rect 219342 3544 219348 3556
rect 219400 3544 219406 3596
rect 236086 3544 236092 3596
rect 236144 3584 236150 3596
rect 237190 3584 237196 3596
rect 236144 3556 237196 3584
rect 236144 3544 236150 3556
rect 237190 3544 237196 3556
rect 237248 3544 237254 3596
rect 237285 3587 237343 3593
rect 237285 3553 237297 3587
rect 237331 3584 237343 3587
rect 293126 3584 293132 3596
rect 237331 3556 293132 3584
rect 237331 3553 237343 3556
rect 237285 3547 237343 3553
rect 293126 3544 293132 3556
rect 293184 3544 293190 3596
rect 304994 3544 305000 3596
rect 305052 3584 305058 3596
rect 306190 3584 306196 3596
rect 305052 3556 306196 3584
rect 305052 3544 305058 3556
rect 306190 3544 306196 3556
rect 306248 3544 306254 3596
rect 310422 3544 310428 3596
rect 310480 3584 310486 3596
rect 365533 3587 365591 3593
rect 365533 3584 365545 3587
rect 310480 3556 365545 3584
rect 310480 3544 310486 3556
rect 365533 3553 365545 3556
rect 365579 3553 365591 3587
rect 365533 3547 365591 3553
rect 365625 3587 365683 3593
rect 365625 3553 365637 3587
rect 365671 3584 365683 3587
rect 368014 3584 368020 3596
rect 365671 3556 368020 3584
rect 365671 3553 365683 3556
rect 365625 3547 365683 3553
rect 368014 3544 368020 3556
rect 368072 3544 368078 3596
rect 415302 3544 415308 3596
rect 415360 3584 415366 3596
rect 475102 3584 475108 3596
rect 415360 3556 475108 3584
rect 415360 3544 415366 3556
rect 475102 3544 475108 3556
rect 475160 3544 475166 3596
rect 494146 3544 494152 3596
rect 494204 3584 494210 3596
rect 495342 3584 495348 3596
rect 494204 3556 495348 3584
rect 494204 3544 494210 3556
rect 495342 3544 495348 3556
rect 495400 3544 495406 3596
rect 517422 3544 517428 3596
rect 517480 3584 517486 3596
rect 577406 3584 577412 3596
rect 517480 3556 577412 3584
rect 517480 3544 517486 3556
rect 577406 3544 577412 3556
rect 577464 3544 577470 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 74350 3476 74356 3528
rect 74408 3516 74414 3528
rect 132497 3519 132555 3525
rect 132497 3516 132509 3519
rect 74408 3488 132509 3516
rect 74408 3476 74414 3488
rect 132497 3485 132509 3488
rect 132543 3485 132555 3519
rect 132497 3479 132555 3485
rect 132586 3476 132592 3528
rect 132644 3516 132650 3528
rect 133782 3516 133788 3528
rect 132644 3488 133788 3516
rect 132644 3476 132650 3488
rect 133782 3476 133788 3488
rect 133840 3476 133846 3528
rect 171042 3476 171048 3528
rect 171100 3516 171106 3528
rect 232498 3516 232504 3528
rect 171100 3488 232504 3516
rect 171100 3476 171106 3488
rect 232498 3476 232504 3488
rect 232556 3476 232562 3528
rect 244274 3476 244280 3528
rect 244332 3516 244338 3528
rect 245562 3516 245568 3528
rect 244332 3488 245568 3516
rect 244332 3476 244338 3488
rect 245562 3476 245568 3488
rect 245620 3476 245626 3528
rect 249702 3476 249708 3528
rect 249760 3516 249766 3528
rect 310974 3516 310980 3528
rect 249760 3488 310980 3516
rect 249760 3476 249766 3488
rect 310974 3476 310980 3488
rect 311032 3476 311038 3528
rect 321462 3476 321468 3528
rect 321520 3516 321526 3528
rect 382366 3516 382372 3528
rect 321520 3488 382372 3516
rect 321520 3476 321526 3488
rect 382366 3476 382372 3488
rect 382424 3476 382430 3528
rect 429102 3476 429108 3528
rect 429160 3516 429166 3528
rect 489362 3516 489368 3528
rect 429160 3488 489368 3516
rect 429160 3476 429166 3488
rect 489362 3476 489368 3488
rect 489420 3476 489426 3528
rect 518802 3476 518808 3528
rect 518860 3516 518866 3528
rect 578602 3516 578608 3528
rect 518860 3488 578608 3516
rect 518860 3476 518866 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 62114 3448 62120 3460
rect 624 3420 62120 3448
rect 624 3408 630 3420
rect 62114 3408 62120 3420
rect 62172 3408 62178 3460
rect 95142 3408 95148 3460
rect 95200 3448 95206 3460
rect 156322 3448 156328 3460
rect 95200 3420 156328 3448
rect 95200 3408 95206 3420
rect 156322 3408 156328 3420
rect 156380 3408 156386 3460
rect 164142 3408 164148 3460
rect 164200 3448 164206 3460
rect 225322 3448 225328 3460
rect 164200 3420 225328 3448
rect 164200 3408 164206 3420
rect 225322 3408 225328 3420
rect 225380 3408 225386 3460
rect 242802 3408 242808 3460
rect 242860 3448 242866 3460
rect 303798 3448 303804 3460
rect 242860 3420 303804 3448
rect 242860 3408 242866 3420
rect 303798 3408 303804 3420
rect 303856 3408 303862 3460
rect 307662 3408 307668 3460
rect 307720 3448 307726 3460
rect 365625 3451 365683 3457
rect 365625 3448 365637 3451
rect 307720 3420 365637 3448
rect 307720 3408 307726 3420
rect 365625 3417 365637 3420
rect 365671 3417 365683 3451
rect 365625 3411 365683 3417
rect 365714 3408 365720 3460
rect 365772 3448 365778 3460
rect 366910 3448 366916 3460
rect 365772 3420 366916 3448
rect 365772 3408 365778 3420
rect 366910 3408 366916 3420
rect 366968 3408 366974 3460
rect 371142 3408 371148 3460
rect 371200 3448 371206 3460
rect 432322 3448 432328 3460
rect 371200 3420 432328 3448
rect 371200 3408 371206 3420
rect 432322 3408 432328 3420
rect 432380 3408 432386 3460
rect 436002 3408 436008 3460
rect 436060 3448 436066 3460
rect 496538 3448 496544 3460
rect 436060 3420 496544 3448
rect 436060 3408 436066 3420
rect 496538 3408 496544 3420
rect 496596 3408 496602 3460
rect 521562 3408 521568 3460
rect 521620 3448 521626 3460
rect 582190 3448 582196 3460
rect 521620 3420 582196 3448
rect 521620 3408 521626 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 125502 3340 125508 3392
rect 125560 3380 125566 3392
rect 183373 3383 183431 3389
rect 183373 3380 183385 3383
rect 125560 3352 183385 3380
rect 125560 3340 125566 3352
rect 183373 3349 183385 3352
rect 183419 3349 183431 3383
rect 183373 3343 183431 3349
rect 183554 3340 183560 3392
rect 183612 3380 183618 3392
rect 184842 3380 184848 3392
rect 183612 3352 184848 3380
rect 183612 3340 183618 3352
rect 184842 3340 184848 3352
rect 184900 3340 184906 3392
rect 204162 3340 204168 3392
rect 204220 3380 204226 3392
rect 264606 3380 264612 3392
rect 204220 3352 264612 3380
rect 204220 3340 204226 3352
rect 264606 3340 264612 3352
rect 264664 3340 264670 3392
rect 270494 3340 270500 3392
rect 270552 3380 270558 3392
rect 271690 3380 271696 3392
rect 270552 3352 271696 3380
rect 270552 3340 270558 3352
rect 271690 3340 271696 3352
rect 271748 3340 271754 3392
rect 287054 3340 287060 3392
rect 287112 3380 287118 3392
rect 288342 3380 288348 3392
rect 287112 3352 288348 3380
rect 287112 3340 287118 3352
rect 288342 3340 288348 3352
rect 288400 3340 288406 3392
rect 293862 3340 293868 3392
rect 293920 3380 293926 3392
rect 353754 3380 353760 3392
rect 293920 3352 353760 3380
rect 293920 3340 293926 3352
rect 353754 3340 353760 3352
rect 353812 3340 353818 3392
rect 357158 3340 357164 3392
rect 357216 3380 357222 3392
rect 417970 3380 417976 3392
rect 357216 3352 417976 3380
rect 357216 3340 357222 3352
rect 417970 3340 417976 3352
rect 418028 3340 418034 3392
rect 451274 3340 451280 3392
rect 451332 3380 451338 3392
rect 452470 3380 452476 3392
rect 451332 3352 452476 3380
rect 451332 3340 451338 3352
rect 452470 3340 452476 3352
rect 452528 3340 452534 3392
rect 467834 3340 467840 3392
rect 467892 3380 467898 3392
rect 469122 3380 469128 3392
rect 467892 3352 469128 3380
rect 467892 3340 467898 3352
rect 469122 3340 469128 3352
rect 469180 3340 469186 3392
rect 471882 3340 471888 3392
rect 471940 3380 471946 3392
rect 532234 3380 532240 3392
rect 471940 3352 532240 3380
rect 471940 3340 471946 3352
rect 532234 3340 532240 3352
rect 532292 3340 532298 3392
rect 536834 3340 536840 3392
rect 536892 3380 536898 3392
rect 538122 3380 538128 3392
rect 536892 3352 538128 3380
rect 536892 3340 536898 3352
rect 538122 3340 538128 3352
rect 538180 3340 538186 3392
rect 571426 3340 571432 3392
rect 571484 3380 571490 3392
rect 572622 3380 572628 3392
rect 571484 3352 572628 3380
rect 571484 3340 571490 3352
rect 572622 3340 572628 3352
rect 572680 3340 572686 3392
rect 132497 3315 132555 3321
rect 132497 3281 132509 3315
rect 132543 3312 132555 3315
rect 136082 3312 136088 3324
rect 132543 3284 136088 3312
rect 132543 3281 132555 3284
rect 132497 3275 132555 3281
rect 136082 3272 136088 3284
rect 136140 3272 136146 3324
rect 136542 3272 136548 3324
rect 136600 3312 136606 3324
rect 196802 3312 196808 3324
rect 136600 3284 196808 3312
rect 136600 3272 136606 3284
rect 196802 3272 196808 3284
rect 196860 3272 196866 3324
rect 215202 3272 215208 3324
rect 215260 3312 215266 3324
rect 275278 3312 275284 3324
rect 215260 3284 275284 3312
rect 215260 3272 215266 3284
rect 275278 3272 275284 3284
rect 275336 3272 275342 3324
rect 343542 3272 343548 3324
rect 343600 3312 343606 3324
rect 403710 3312 403716 3324
rect 343600 3284 403716 3312
rect 343600 3272 343606 3284
rect 403710 3272 403716 3284
rect 403768 3272 403774 3324
rect 478782 3272 478788 3324
rect 478840 3312 478846 3324
rect 539318 3312 539324 3324
rect 478840 3284 539324 3312
rect 478840 3272 478846 3284
rect 539318 3272 539324 3284
rect 539376 3272 539382 3324
rect 100662 3204 100668 3256
rect 100720 3244 100726 3256
rect 161106 3244 161112 3256
rect 100720 3216 161112 3244
rect 100720 3204 100726 3216
rect 161106 3204 161112 3216
rect 161164 3204 161170 3256
rect 175366 3204 175372 3256
rect 175424 3244 175430 3256
rect 176562 3244 176568 3256
rect 175424 3216 176568 3244
rect 175424 3204 175430 3216
rect 176562 3204 176568 3216
rect 176620 3204 176626 3256
rect 183373 3247 183431 3253
rect 183373 3213 183385 3247
rect 183419 3244 183431 3247
rect 186038 3244 186044 3256
rect 183419 3216 186044 3244
rect 183419 3213 183431 3216
rect 183373 3207 183431 3213
rect 186038 3204 186044 3216
rect 186096 3204 186102 3256
rect 193122 3204 193128 3256
rect 193180 3244 193186 3256
rect 253842 3244 253848 3256
rect 193180 3216 253848 3244
rect 193180 3204 193186 3216
rect 253842 3204 253848 3216
rect 253900 3204 253906 3256
rect 314654 3204 314660 3256
rect 314712 3244 314718 3256
rect 375190 3244 375196 3256
rect 314712 3216 375196 3244
rect 314712 3204 314718 3216
rect 375190 3204 375196 3216
rect 375248 3204 375254 3256
rect 460842 3204 460848 3256
rect 460900 3244 460906 3256
rect 521470 3244 521476 3256
rect 460900 3216 521476 3244
rect 460900 3204 460906 3216
rect 521470 3204 521476 3216
rect 521528 3204 521534 3256
rect 107562 3136 107568 3188
rect 107620 3176 107626 3188
rect 168190 3176 168196 3188
rect 107620 3148 168196 3176
rect 107620 3136 107626 3148
rect 168190 3136 168196 3148
rect 168248 3136 168254 3188
rect 186222 3136 186228 3188
rect 186280 3176 186286 3188
rect 246758 3176 246764 3188
rect 186280 3148 246764 3176
rect 186280 3136 186286 3148
rect 246758 3136 246764 3148
rect 246816 3136 246822 3188
rect 332502 3136 332508 3188
rect 332560 3176 332566 3188
rect 393038 3176 393044 3188
rect 332560 3148 393044 3176
rect 332560 3136 332566 3148
rect 393038 3136 393044 3148
rect 393096 3136 393102 3188
rect 453942 3136 453948 3188
rect 454000 3176 454006 3188
rect 514386 3176 514392 3188
rect 454000 3148 514392 3176
rect 454000 3136 454006 3148
rect 514386 3136 514392 3148
rect 514444 3136 514450 3188
rect 92382 3068 92388 3120
rect 92440 3108 92446 3120
rect 152734 3108 152740 3120
rect 92440 3080 152740 3108
rect 92440 3068 92446 3080
rect 152734 3068 152740 3080
rect 152792 3068 152798 3120
rect 222102 3068 222108 3120
rect 222160 3108 222166 3120
rect 282454 3108 282460 3120
rect 222160 3080 282460 3108
rect 222160 3068 222166 3080
rect 282454 3068 282460 3080
rect 282512 3068 282518 3120
rect 336642 3068 336648 3120
rect 336700 3108 336706 3120
rect 396626 3108 396632 3120
rect 336700 3080 396632 3108
rect 336700 3068 336706 3080
rect 396626 3068 396632 3080
rect 396684 3068 396690 3120
rect 458082 3068 458088 3120
rect 458140 3108 458146 3120
rect 517882 3108 517888 3120
rect 458140 3080 517888 3108
rect 458140 3068 458146 3080
rect 517882 3068 517888 3080
rect 517940 3068 517946 3120
rect 99282 3000 99288 3052
rect 99340 3040 99346 3052
rect 159910 3040 159916 3052
rect 99340 3012 159916 3040
rect 99340 3000 99346 3012
rect 159910 3000 159916 3012
rect 159968 3000 159974 3052
rect 365533 3043 365591 3049
rect 365533 3009 365545 3043
rect 365579 3040 365591 3043
rect 371602 3040 371608 3052
rect 365579 3012 371608 3040
rect 365579 3009 365591 3012
rect 365533 3003 365591 3009
rect 371602 3000 371608 3012
rect 371660 3000 371666 3052
rect 464982 3000 464988 3052
rect 465040 3040 465046 3052
rect 525058 3040 525064 3052
rect 465040 3012 525064 3040
rect 465040 3000 465046 3012
rect 525058 3000 525064 3012
rect 525116 3000 525122 3052
rect 440142 2932 440148 2984
rect 440200 2972 440206 2984
rect 500126 2972 500132 2984
rect 440200 2944 500132 2972
rect 440200 2932 440206 2944
rect 500126 2932 500132 2944
rect 500184 2932 500190 2984
rect 433150 2864 433156 2916
rect 433208 2904 433214 2916
rect 492950 2904 492956 2916
rect 433208 2876 492956 2904
rect 433208 2864 433214 2876
rect 492950 2864 492956 2876
rect 493008 2864 493014 2916
rect 393314 2796 393320 2848
rect 393372 2836 393378 2848
rect 393372 2808 394280 2836
rect 393372 2796 393378 2808
rect 394252 2780 394280 2808
rect 394694 2796 394700 2848
rect 394752 2836 394758 2848
rect 394752 2808 395476 2836
rect 394752 2796 394758 2808
rect 395448 2780 395476 2808
rect 397454 2796 397460 2848
rect 397512 2836 397518 2848
rect 397512 2808 397868 2836
rect 397512 2796 397518 2808
rect 397840 2780 397868 2808
rect 412634 2796 412640 2848
rect 412692 2836 412698 2848
rect 412692 2808 413324 2836
rect 412692 2796 412698 2808
rect 413296 2780 413324 2808
rect 419534 2796 419540 2848
rect 419592 2836 419598 2848
rect 419592 2808 420408 2836
rect 419592 2796 419598 2808
rect 420380 2780 420408 2808
rect 426434 2796 426440 2848
rect 426492 2836 426498 2848
rect 426492 2808 427584 2836
rect 426492 2796 426498 2808
rect 427556 2780 427584 2808
rect 427906 2796 427912 2848
rect 427964 2836 427970 2848
rect 427964 2808 428780 2836
rect 427964 2796 427970 2808
rect 428752 2780 428780 2808
rect 430574 2796 430580 2848
rect 430632 2836 430638 2848
rect 430632 2808 431172 2836
rect 430632 2796 430638 2808
rect 431144 2780 431172 2808
rect 394234 2728 394240 2780
rect 394292 2728 394298 2780
rect 395430 2728 395436 2780
rect 395488 2728 395494 2780
rect 397822 2728 397828 2780
rect 397880 2728 397886 2780
rect 413278 2728 413284 2780
rect 413336 2728 413342 2780
rect 420362 2728 420368 2780
rect 420420 2728 420426 2780
rect 427538 2728 427544 2780
rect 427596 2728 427602 2780
rect 428734 2728 428740 2780
rect 428792 2728 428798 2780
rect 431126 2728 431132 2780
rect 431184 2728 431190 2780
rect 347774 2048 347780 2100
rect 347832 2088 347838 2100
rect 349062 2088 349068 2100
rect 347832 2060 349068 2088
rect 347832 2048 347838 2060
rect 349062 2048 349068 2060
rect 349120 2048 349126 2100
rect 375374 552 375380 604
rect 375432 592 375438 604
rect 376386 592 376392 604
rect 375432 564 376392 592
rect 375432 552 375438 564
rect 376386 552 376392 564
rect 376444 552 376450 604
rect 376754 552 376760 604
rect 376812 592 376818 604
rect 377582 592 377588 604
rect 376812 564 377588 592
rect 376812 552 376818 564
rect 377582 552 377588 564
rect 377640 552 377646 604
rect 383654 552 383660 604
rect 383712 592 383718 604
rect 384666 592 384672 604
rect 383712 564 384672 592
rect 383712 552 383718 564
rect 384666 552 384672 564
rect 384724 552 384730 604
rect 386414 552 386420 604
rect 386472 592 386478 604
rect 387058 592 387064 604
rect 386472 564 387064 592
rect 386472 552 386478 564
rect 387058 552 387064 564
rect 387116 552 387122 604
rect 387794 552 387800 604
rect 387852 592 387858 604
rect 388254 592 388260 604
rect 387852 564 388260 592
rect 387852 552 387858 564
rect 388254 552 388260 564
rect 388312 552 388318 604
rect 405734 552 405740 604
rect 405792 592 405798 604
rect 406102 592 406108 604
rect 405792 564 406108 592
rect 405792 552 405798 564
rect 406102 552 406108 564
rect 406160 552 406166 604
rect 412082 592 412088 604
rect 412043 564 412088 592
rect 412082 552 412088 564
rect 412140 552 412146 604
rect 415670 592 415676 604
rect 415631 564 415676 592
rect 415670 552 415676 564
rect 415728 552 415734 604
rect 435818 592 435824 604
rect 435779 564 435824 592
rect 435818 552 435824 564
rect 435876 552 435882 604
rect 455414 552 455420 604
rect 455472 592 455478 604
rect 456058 592 456064 604
rect 455472 564 456064 592
rect 455472 552 455478 564
rect 456058 552 456064 564
rect 456116 552 456122 604
rect 456886 552 456892 604
rect 456944 592 456950 604
rect 457254 592 457260 604
rect 456944 564 457260 592
rect 456944 552 456950 564
rect 457254 552 457260 564
rect 457312 552 457318 604
rect 471974 552 471980 604
rect 472032 592 472038 604
rect 472710 592 472716 604
rect 472032 564 472716 592
rect 472032 552 472038 564
rect 472710 552 472716 564
rect 472768 552 472774 604
rect 473354 552 473360 604
rect 473412 592 473418 604
rect 473906 592 473912 604
rect 473412 564 473912 592
rect 473412 552 473418 564
rect 473906 552 473912 564
rect 473964 552 473970 604
rect 478874 552 478880 604
rect 478932 592 478938 604
rect 479886 592 479892 604
rect 478932 564 479892 592
rect 478932 552 478938 564
rect 479886 552 479892 564
rect 479944 552 479950 604
rect 579614 552 579620 604
rect 579672 592 579678 604
rect 579798 592 579804 604
rect 579672 564 579804 592
rect 579672 552 579678 564
rect 579798 552 579804 564
rect 579856 552 579862 604
<< via1 >>
rect 394608 700408 394660 700460
rect 413652 700408 413704 700460
rect 463608 700408 463660 700460
rect 494796 700408 494848 700460
rect 514668 700408 514720 700460
rect 559656 700408 559708 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 411168 700340 411220 700392
rect 429844 700340 429896 700392
rect 445668 700340 445720 700392
rect 478512 700340 478564 700392
rect 496728 700340 496780 700392
rect 543464 700340 543516 700392
rect 344284 700272 344336 700324
rect 348792 700272 348844 700324
rect 378048 700272 378100 700324
rect 397460 700272 397512 700324
rect 429108 700272 429160 700324
rect 462320 700272 462372 700324
rect 480168 700272 480220 700324
rect 527180 700272 527232 700324
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 326988 699660 327040 699712
rect 332508 699660 332560 699712
rect 360108 699660 360160 699712
rect 364984 699660 365036 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 137744 698232 137796 698284
rect 137928 698232 137980 698284
rect 523776 696940 523828 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 283840 695512 283892 695564
rect 283932 695512 283984 695564
rect 8208 695444 8260 695496
rect 137928 695444 137980 695496
rect 219164 695444 219216 695496
rect 72700 694084 72752 694136
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 283932 688576 283984 688628
rect 284116 688576 284168 688628
rect 8116 685899 8168 685908
rect 8116 685865 8125 685899
rect 8125 685865 8159 685899
rect 8159 685865 8168 685899
rect 8116 685856 8168 685865
rect 137836 685899 137888 685908
rect 137836 685865 137845 685899
rect 137845 685865 137879 685899
rect 137879 685865 137888 685899
rect 137836 685856 137888 685865
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 523684 685856 523736 685908
rect 580172 685856 580224 685908
rect 154396 685788 154448 685840
rect 284116 685788 284168 685840
rect 72516 684607 72568 684616
rect 72516 684573 72525 684607
rect 72525 684573 72559 684607
rect 72559 684573 72568 684607
rect 72516 684564 72568 684573
rect 72516 684428 72568 684480
rect 8116 678988 8168 679040
rect 137836 678988 137888 679040
rect 8024 678920 8076 678972
rect 137744 678920 137796 678972
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 284024 676243 284076 676252
rect 284024 676209 284033 676243
rect 284033 676209 284067 676243
rect 284067 676209 284076 676243
rect 284024 676200 284076 676209
rect 218980 676175 219032 676184
rect 218980 676141 218989 676175
rect 218989 676141 219023 676175
rect 219023 676141 219032 676175
rect 218980 676132 219032 676141
rect 72792 676107 72844 676116
rect 72792 676073 72801 676107
rect 72801 676073 72835 676107
rect 72835 676073 72844 676107
rect 72792 676064 72844 676073
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 137744 673480 137796 673532
rect 137928 673480 137980 673532
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 284024 673480 284076 673532
rect 284208 673480 284260 673532
rect 72792 669332 72844 669384
rect 72792 669196 72844 669248
rect 219072 666544 219124 666596
rect 8024 654100 8076 654152
rect 8208 654100 8260 654152
rect 137744 654100 137796 654152
rect 137928 654100 137980 654152
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 284024 654100 284076 654152
rect 284208 654100 284260 654152
rect 342996 645804 343048 645856
rect 344284 645804 344336 645856
rect 377128 645804 377180 645856
rect 378048 645804 378100 645856
rect 428188 645804 428240 645856
rect 429108 645804 429160 645856
rect 462320 645804 462372 645856
rect 463608 645804 463660 645856
rect 479340 645804 479392 645856
rect 480168 645804 480220 645856
rect 513380 645600 513432 645652
rect 514668 645600 514720 645652
rect 325976 645464 326028 645516
rect 326988 645464 327040 645516
rect 73068 645328 73120 645380
rect 121552 645328 121604 645380
rect 137928 645328 137980 645380
rect 172704 645328 172756 645380
rect 8208 645260 8260 645312
rect 70492 645260 70544 645312
rect 89628 645260 89680 645312
rect 138572 645260 138624 645312
rect 41328 645192 41380 645244
rect 104532 645192 104584 645244
rect 154488 645192 154540 645244
rect 189724 645192 189776 645244
rect 202788 645192 202840 645244
rect 223764 645192 223816 645244
rect 235908 645192 235960 645244
rect 257896 645192 257948 645244
rect 24768 645124 24820 645176
rect 87512 645124 87564 645176
rect 106188 645124 106240 645176
rect 155592 645124 155644 645176
rect 171048 645124 171100 645176
rect 206744 645124 206796 645176
rect 219348 645124 219400 645176
rect 240784 645124 240836 645176
rect 267648 645124 267700 645176
rect 274916 645124 274968 645176
rect 284208 645124 284260 645176
rect 291936 645124 291988 645176
rect 300768 644852 300820 644904
rect 308956 644852 309008 644904
rect 523868 638936 523920 638988
rect 580172 638936 580224 638988
rect 3424 636148 3476 636200
rect 59360 636148 59412 636200
rect 3516 622344 3568 622396
rect 59360 622344 59412 622396
rect 524328 609900 524380 609952
rect 580264 609900 580316 609952
rect 3608 608540 3660 608592
rect 59360 608540 59412 608592
rect 523776 603100 523828 603152
rect 580172 603100 580224 603152
rect 523684 597456 523736 597508
rect 580448 597456 580500 597508
rect 3424 593308 3476 593360
rect 59360 593308 59412 593360
rect 523684 592016 523736 592068
rect 580172 592016 580224 592068
rect 3516 579572 3568 579624
rect 59360 579572 59412 579624
rect 524328 569848 524380 569900
rect 580356 569848 580408 569900
rect 3608 565768 3660 565820
rect 59360 565768 59412 565820
rect 523868 556180 523920 556232
rect 580172 556180 580224 556232
rect 3424 550536 3476 550588
rect 59360 550536 59412 550588
rect 523776 545096 523828 545148
rect 580172 545096 580224 545148
rect 3516 536732 3568 536784
rect 59360 536732 59412 536784
rect 523224 531224 523276 531276
rect 580264 531224 580316 531276
rect 3424 522928 3476 522980
rect 59360 522928 59412 522980
rect 523868 509260 523920 509312
rect 580172 509260 580224 509312
rect 3332 507764 3384 507816
rect 59360 507764 59412 507816
rect 523776 498176 523828 498228
rect 580172 498176 580224 498228
rect 3332 493960 3384 494012
rect 59360 493960 59412 494012
rect 524328 491240 524380 491292
rect 580356 491240 580408 491292
rect 523684 485800 523736 485852
rect 580172 485800 580224 485852
rect 3608 480156 3660 480208
rect 59360 480156 59412 480208
rect 3424 463700 3476 463752
rect 59360 463700 59412 463752
rect 523868 462340 523920 462392
rect 580172 462340 580224 462392
rect 523776 451256 523828 451308
rect 580172 451256 580224 451308
rect 3424 449896 3476 449948
rect 59360 449896 59412 449948
rect 523684 438880 523736 438932
rect 580172 438880 580224 438932
rect 3424 436092 3476 436144
rect 59360 436092 59412 436144
rect 3516 420928 3568 420980
rect 59360 420928 59412 420980
rect 523868 415420 523920 415472
rect 580172 415420 580224 415472
rect 3424 407124 3476 407176
rect 59360 407124 59412 407176
rect 523776 404336 523828 404388
rect 580172 404336 580224 404388
rect 3516 391960 3568 392012
rect 59360 391960 59412 392012
rect 523684 391960 523736 392012
rect 580172 391960 580224 392012
rect 3424 378156 3476 378208
rect 59360 378156 59412 378208
rect 523684 368500 523736 368552
rect 580172 368500 580224 368552
rect 3516 364352 3568 364404
rect 59360 364352 59412 364404
rect 523776 357416 523828 357468
rect 580172 357416 580224 357468
rect 3608 349120 3660 349172
rect 59360 349120 59412 349172
rect 523684 345040 523736 345092
rect 580172 345040 580224 345092
rect 3424 335316 3476 335368
rect 59360 335316 59412 335368
rect 3516 321580 3568 321632
rect 59360 321580 59412 321632
rect 523500 321580 523552 321632
rect 580172 321580 580224 321632
rect 523684 310496 523736 310548
rect 579804 310496 579856 310548
rect 3700 306348 3752 306400
rect 59360 306348 59412 306400
rect 523224 298120 523276 298172
rect 580172 298120 580224 298172
rect 3608 292544 3660 292596
rect 59360 292544 59412 292596
rect 3424 278740 3476 278792
rect 59360 278740 59412 278792
rect 524328 275952 524380 276004
rect 580172 275952 580224 276004
rect 3700 263576 3752 263628
rect 59360 263576 59412 263628
rect 524328 263576 524380 263628
rect 579804 263576 579856 263628
rect 523960 251200 524012 251252
rect 580172 251200 580224 251252
rect 3516 249772 3568 249824
rect 59360 249772 59412 249824
rect 3608 235968 3660 236020
rect 59360 235968 59412 236020
rect 523684 229032 523736 229084
rect 580172 229032 580224 229084
rect 3424 220804 3476 220856
rect 59360 220804 59412 220856
rect 523684 217948 523736 218000
rect 580172 217948 580224 218000
rect 3700 207000 3752 207052
rect 59360 207000 59412 207052
rect 523408 205572 523460 205624
rect 579804 205572 579856 205624
rect 3608 191836 3660 191888
rect 59360 191836 59412 191888
rect 523684 182112 523736 182164
rect 580172 182112 580224 182164
rect 3516 178032 3568 178084
rect 59360 178032 59412 178084
rect 523776 171028 523828 171080
rect 580172 171028 580224 171080
rect 3424 164228 3476 164280
rect 59360 164228 59412 164280
rect 523684 158652 523736 158704
rect 579804 158652 579856 158704
rect 3700 149064 3752 149116
rect 59360 149064 59412 149116
rect 3608 135260 3660 135312
rect 59360 135260 59412 135312
rect 523684 135192 523736 135244
rect 580172 135192 580224 135244
rect 523868 124108 523920 124160
rect 580172 124108 580224 124160
rect 3516 121456 3568 121508
rect 59360 121456 59412 121508
rect 523776 111732 523828 111784
rect 579804 111732 579856 111784
rect 3792 106292 3844 106344
rect 59360 106292 59412 106344
rect 3700 92488 3752 92540
rect 59360 92488 59412 92540
rect 523684 88272 523736 88324
rect 580172 88272 580224 88324
rect 3424 78684 3476 78736
rect 59360 78684 59412 78736
rect 523776 77188 523828 77240
rect 580172 77188 580224 77240
rect 523868 64812 523920 64864
rect 579804 64812 579856 64864
rect 3608 63520 3660 63572
rect 59360 63520 59412 63572
rect 3516 49716 3568 49768
rect 59360 49716 59412 49768
rect 523684 41352 523736 41404
rect 580172 41352 580224 41404
rect 272248 41216 272300 41268
rect 273168 41216 273220 41268
rect 369952 41216 370004 41268
rect 371056 41216 371108 41268
rect 145932 41148 145984 41200
rect 167368 41148 167420 41200
rect 227904 41148 227956 41200
rect 253204 41148 253256 41200
rect 110236 41080 110288 41132
rect 171232 41080 171284 41132
rect 188896 41080 188948 41132
rect 249892 41080 249944 41132
rect 396172 41080 396224 41132
rect 456892 41080 456944 41132
rect 131672 41012 131724 41064
rect 193404 41012 193456 41064
rect 81624 40944 81676 40996
rect 142252 40944 142304 40996
rect 207112 40944 207164 40996
rect 210332 40944 210384 40996
rect 270500 40944 270552 40996
rect 318708 41012 318760 41064
rect 343732 41012 343784 41064
rect 344836 41012 344888 41064
rect 367652 41012 367704 41064
rect 403348 41012 403400 41064
rect 463792 41012 463844 41064
rect 427912 40944 427964 40996
rect 103060 40876 103112 40928
rect 164332 40876 164384 40928
rect 174544 40876 174596 40928
rect 236184 40876 236236 40928
rect 267648 40876 267700 40928
rect 328552 40876 328604 40928
rect 345664 40876 345716 40928
rect 374736 40876 374788 40928
rect 434812 40876 434864 40928
rect 474832 40876 474884 40928
rect 535460 40876 535512 40928
rect 95884 40808 95936 40860
rect 157432 40808 157484 40860
rect 181720 40808 181772 40860
rect 242992 40808 243044 40860
rect 260380 40808 260432 40860
rect 321744 40808 321796 40860
rect 381912 40808 381964 40860
rect 443184 40808 443236 40860
rect 489184 40808 489236 40860
rect 549260 40808 549312 40860
rect 88708 40740 88760 40792
rect 150624 40740 150676 40792
rect 224592 40740 224644 40792
rect 285772 40740 285824 40792
rect 333060 40740 333112 40792
rect 333888 40740 333940 40792
rect 334256 40740 334308 40792
rect 367744 40740 367796 40792
rect 389088 40740 389140 40792
rect 449992 40740 450044 40792
rect 459376 40740 459428 40792
rect 467104 40740 467156 40792
rect 482008 40740 482060 40792
rect 542360 40740 542412 40792
rect 2688 40672 2740 40724
rect 63684 40672 63736 40724
rect 67272 40672 67324 40724
rect 128452 40672 128504 40724
rect 138848 40672 138900 40724
rect 200212 40672 200264 40724
rect 217416 40672 217468 40724
rect 278964 40672 279016 40724
rect 316408 40672 316460 40724
rect 317328 40672 317380 40724
rect 324688 40672 324740 40724
rect 325608 40672 325660 40724
rect 346124 40672 346176 40724
rect 407212 40672 407264 40724
rect 467748 40672 467800 40724
rect 528560 40672 528612 40724
rect 378324 40604 378376 40656
rect 379428 40604 379480 40656
rect 247224 40536 247276 40588
rect 248328 40536 248380 40588
rect 299664 40536 299716 40588
rect 300768 40536 300820 40588
rect 290188 40468 290240 40520
rect 291108 40468 291160 40520
rect 300860 40468 300912 40520
rect 302148 40468 302200 40520
rect 283012 40332 283064 40384
rect 284208 40332 284260 40384
rect 313464 40332 313516 40384
rect 335452 40332 335504 40384
rect 336648 40332 336700 40384
rect 64880 40128 64932 40180
rect 66168 40128 66220 40180
rect 66076 40060 66128 40112
rect 66904 40060 66956 40112
rect 70860 40060 70912 40112
rect 71688 40060 71740 40112
rect 72056 40060 72108 40112
rect 73068 40060 73120 40112
rect 80428 40060 80480 40112
rect 81348 40060 81400 40112
rect 82820 40060 82872 40112
rect 84016 40060 84068 40112
rect 89904 40060 89956 40112
rect 91008 40060 91060 40112
rect 91100 40060 91152 40112
rect 92388 40060 92440 40112
rect 97080 40060 97132 40112
rect 97908 40060 97960 40112
rect 98276 40060 98328 40112
rect 99288 40060 99340 40112
rect 99472 40060 99524 40112
rect 100668 40060 100720 40112
rect 105452 40060 105504 40112
rect 106188 40060 106240 40112
rect 106648 40060 106700 40112
rect 107568 40060 107620 40112
rect 107844 40060 107896 40112
rect 108948 40060 109000 40112
rect 109040 40060 109092 40112
rect 110328 40060 110380 40112
rect 113732 40060 113784 40112
rect 114468 40060 114520 40112
rect 114928 40060 114980 40112
rect 115848 40060 115900 40112
rect 116124 40060 116176 40112
rect 117228 40060 117280 40112
rect 117320 40060 117372 40112
rect 118608 40060 118660 40112
rect 124496 40060 124548 40112
rect 125508 40060 125560 40112
rect 125692 40060 125744 40112
rect 126796 40060 126848 40112
rect 132868 40060 132920 40112
rect 133788 40060 133840 40112
rect 134064 40060 134116 40112
rect 135168 40060 135220 40112
rect 135260 40060 135312 40112
rect 136548 40060 136600 40112
rect 141148 40060 141200 40112
rect 142068 40060 142120 40112
rect 142344 40060 142396 40112
rect 143448 40060 143500 40112
rect 143540 40060 143592 40112
rect 144828 40060 144880 40112
rect 149520 40060 149572 40112
rect 150348 40060 150400 40112
rect 150716 40060 150768 40112
rect 151728 40060 151780 40112
rect 157892 40060 157944 40112
rect 158628 40060 158680 40112
rect 160284 40060 160336 40112
rect 161388 40060 161440 40112
rect 161480 40060 161532 40112
rect 162768 40060 162820 40112
rect 166172 40060 166224 40112
rect 166908 40060 166960 40112
rect 168564 40060 168616 40112
rect 169668 40060 169720 40112
rect 169760 40060 169812 40112
rect 170956 40060 171008 40112
rect 175740 40060 175792 40112
rect 176568 40060 176620 40112
rect 176936 40060 176988 40112
rect 177948 40060 178000 40112
rect 178132 40060 178184 40112
rect 179328 40060 179380 40112
rect 185308 40060 185360 40112
rect 186228 40060 186280 40112
rect 186504 40060 186556 40112
rect 187608 40060 187660 40112
rect 193588 40060 193640 40112
rect 194508 40060 194560 40112
rect 195980 40060 196032 40112
rect 197268 40060 197320 40112
rect 201960 40060 202012 40112
rect 202788 40060 202840 40112
rect 203156 40060 203208 40112
rect 204168 40060 204220 40112
rect 204352 40060 204404 40112
rect 205548 40060 205600 40112
rect 211528 40060 211580 40112
rect 212448 40060 212500 40112
rect 212724 40060 212776 40112
rect 213828 40060 213880 40112
rect 213920 40060 213972 40112
rect 215208 40060 215260 40112
rect 218612 40060 218664 40112
rect 219348 40060 219400 40112
rect 221004 40060 221056 40112
rect 222108 40060 222160 40112
rect 222200 40060 222252 40112
rect 223488 40060 223540 40112
rect 228180 40060 228232 40112
rect 229008 40060 229060 40112
rect 229376 40060 229428 40112
rect 230388 40060 230440 40112
rect 230572 40060 230624 40112
rect 231676 40060 231728 40112
rect 237748 40060 237800 40112
rect 238668 40060 238720 40112
rect 238944 40060 238996 40112
rect 240048 40060 240100 40112
rect 240140 40060 240192 40112
rect 241428 40060 241480 40112
rect 246028 40060 246080 40112
rect 246948 40060 247000 40112
rect 254400 40060 254452 40112
rect 255228 40060 255280 40112
rect 255596 40060 255648 40112
rect 256608 40060 256660 40112
rect 256792 40060 256844 40112
rect 257988 40060 258040 40112
rect 262772 40060 262824 40112
rect 263508 40060 263560 40112
rect 263968 40060 264020 40112
rect 264888 40060 264940 40112
rect 265164 40060 265216 40112
rect 266268 40060 266320 40112
rect 271052 40060 271104 40112
rect 272524 40060 272576 40112
rect 274640 40060 274692 40112
rect 275836 40060 275888 40112
rect 281816 40060 281868 40112
rect 282828 40060 282880 40112
rect 291384 40060 291436 40112
rect 292488 40060 292540 40112
rect 292580 40060 292632 40112
rect 293868 40060 293920 40112
rect 306840 40060 306892 40112
rect 307668 40060 307720 40112
rect 308036 40060 308088 40112
rect 309048 40060 309100 40112
rect 309232 40060 309284 40112
rect 311164 40060 311216 40112
rect 315212 40060 315264 40112
rect 315948 40060 316000 40112
rect 317604 40060 317656 40112
rect 318708 40060 318760 40112
rect 323492 40060 323544 40112
rect 324228 40060 324280 40112
rect 325884 40060 325936 40112
rect 326988 40060 327040 40112
rect 342628 40060 342680 40112
rect 343548 40060 343600 40112
rect 350908 40060 350960 40112
rect 351828 40060 351880 40112
rect 352104 40060 352156 40112
rect 353208 40060 353260 40112
rect 353300 40060 353352 40112
rect 354588 40060 354640 40112
rect 360476 40060 360528 40112
rect 361488 40060 361540 40112
rect 361672 40060 361724 40112
rect 362868 40060 362920 40112
rect 368848 40060 368900 40112
rect 369768 40060 369820 40112
rect 375932 40060 375984 40112
rect 376668 40060 376720 40112
rect 377128 40060 377180 40112
rect 378048 40060 378100 40112
rect 379520 40060 379572 40112
rect 380808 40060 380860 40112
rect 385500 40060 385552 40112
rect 386328 40060 386380 40112
rect 386696 40060 386748 40112
rect 387708 40060 387760 40112
rect 387892 40060 387944 40112
rect 389088 40060 389140 40112
rect 394976 40060 395028 40112
rect 395988 40060 396040 40112
rect 404544 40060 404596 40112
rect 405648 40060 405700 40112
rect 405740 40060 405792 40112
rect 406936 40060 406988 40112
rect 411720 40060 411772 40112
rect 412548 40060 412600 40112
rect 412916 40060 412968 40112
rect 413928 40060 413980 40112
rect 414112 40060 414164 40112
rect 415308 40060 415360 40112
rect 420092 40060 420144 40112
rect 420828 40060 420880 40112
rect 421196 40060 421248 40112
rect 422208 40060 422260 40112
rect 422392 40060 422444 40112
rect 423588 40060 423640 40112
rect 428372 40060 428424 40112
rect 429108 40060 429160 40112
rect 429568 40060 429620 40112
rect 430488 40060 430540 40112
rect 430764 40060 430816 40112
rect 431868 40060 431920 40112
rect 431960 40060 432012 40112
rect 433156 40060 433208 40112
rect 437940 40060 437992 40112
rect 438768 40060 438820 40112
rect 439136 40060 439188 40112
rect 440148 40060 440200 40112
rect 440332 40060 440384 40112
rect 441528 40060 441580 40112
rect 446220 40060 446272 40112
rect 447048 40060 447100 40112
rect 447416 40060 447468 40112
rect 448428 40060 448480 40112
rect 448612 40060 448664 40112
rect 449716 40060 449768 40112
rect 455788 40060 455840 40112
rect 456708 40060 456760 40112
rect 456984 40060 457036 40112
rect 458088 40060 458140 40112
rect 458180 40060 458232 40112
rect 459468 40060 459520 40112
rect 464160 40060 464212 40112
rect 464988 40060 465040 40112
rect 465356 40060 465408 40112
rect 466368 40060 466420 40112
rect 466552 40060 466604 40112
rect 467748 40060 467800 40112
rect 472440 40060 472492 40112
rect 473268 40060 473320 40112
rect 473636 40060 473688 40112
rect 474648 40060 474700 40112
rect 480812 40060 480864 40112
rect 481548 40060 481600 40112
rect 483204 40060 483256 40112
rect 484308 40060 484360 40112
rect 484400 40060 484452 40112
rect 485596 40060 485648 40112
rect 490380 40060 490432 40112
rect 491208 40060 491260 40112
rect 491576 40060 491628 40112
rect 492588 40060 492640 40112
rect 492772 40060 492824 40112
rect 493968 40060 494020 40112
rect 498660 40060 498712 40112
rect 499488 40060 499540 40112
rect 499856 40060 499908 40112
rect 500868 40060 500920 40112
rect 508228 40060 508280 40112
rect 509148 40060 509200 40112
rect 509424 40060 509476 40112
rect 510528 40060 510580 40112
rect 510620 40060 510672 40112
rect 511908 40060 511960 40112
rect 516600 40060 516652 40112
rect 517428 40060 517480 40112
rect 517796 40060 517848 40112
rect 518808 40060 518860 40112
rect 287796 39448 287848 39500
rect 347780 39448 347832 39500
rect 73252 39380 73304 39432
rect 133880 39380 133932 39432
rect 159088 39380 159140 39432
rect 219440 39380 219492 39432
rect 226984 39380 227036 39432
rect 287060 39380 287112 39432
rect 319904 39380 319956 39432
rect 380900 39380 380952 39432
rect 126888 39312 126940 39364
rect 187700 39312 187752 39364
rect 194784 39312 194836 39364
rect 255320 39312 255372 39364
rect 259184 39312 259236 39364
rect 320180 39312 320232 39364
rect 366456 39312 366508 39364
rect 426440 39312 426492 39364
rect 433248 39312 433300 39364
rect 494060 39312 494112 39364
rect 501052 39312 501104 39364
rect 561680 39312 561732 39364
rect 434812 38607 434864 38616
rect 434812 38573 434821 38607
rect 434821 38573 434855 38607
rect 434855 38573 434864 38607
rect 434812 38564 434864 38573
rect 187976 38020 188028 38072
rect 248420 38020 248472 38072
rect 402152 38020 402204 38072
rect 462320 38020 462372 38072
rect 123300 37952 123352 38004
rect 183560 37952 183612 38004
rect 219808 37952 219860 38004
rect 280160 37952 280212 38004
rect 280620 37952 280672 38004
rect 340880 37952 340932 38004
rect 359280 37952 359332 38004
rect 419540 37952 419592 38004
rect 76840 37884 76892 37936
rect 138020 37884 138072 37936
rect 155500 37884 155552 37936
rect 216680 37884 216732 37936
rect 248696 37884 248748 37936
rect 309140 37884 309192 37936
rect 312820 37884 312872 37936
rect 374092 37884 374144 37936
rect 451004 37884 451056 37936
rect 512000 37884 512052 37936
rect 518992 37884 519044 37936
rect 579620 37884 579672 37936
rect 184112 36660 184164 36712
rect 244280 36660 244332 36712
rect 244832 36660 244884 36712
rect 305000 36660 305052 36712
rect 305644 36660 305696 36712
rect 365720 36660 365772 36712
rect 151912 36592 151964 36644
rect 212540 36592 212592 36644
rect 277032 36592 277084 36644
rect 338120 36592 338172 36644
rect 119712 36524 119764 36576
rect 180800 36524 180852 36576
rect 216220 36524 216272 36576
rect 277400 36524 277452 36576
rect 348516 36524 348568 36576
rect 408500 36524 408552 36576
rect 415216 36524 415268 36576
rect 476120 36524 476172 36576
rect 493876 36524 493928 36576
rect 554780 36524 554832 36576
rect 213828 35300 213880 35352
rect 273260 35300 273312 35352
rect 273444 35300 273496 35352
rect 333980 35300 334032 35352
rect 117228 35232 117280 35284
rect 176660 35232 176712 35284
rect 180708 35232 180760 35284
rect 241520 35232 241572 35284
rect 302056 35232 302108 35284
rect 362960 35232 363012 35284
rect 391848 35232 391900 35284
rect 451280 35232 451332 35284
rect 148968 35164 149020 35216
rect 209872 35164 209924 35216
rect 241336 35164 241388 35216
rect 302240 35164 302292 35216
rect 342168 35164 342220 35216
rect 401600 35164 401652 35216
rect 413928 35164 413980 35216
rect 473360 35164 473412 35216
rect 511816 35164 511868 35216
rect 571432 35164 571484 35216
rect 177948 33872 178000 33924
rect 237380 33872 237432 33924
rect 238668 33872 238720 33924
rect 298100 33872 298152 33924
rect 113088 33804 113140 33856
rect 173900 33804 173952 33856
rect 205456 33804 205508 33856
rect 266360 33804 266412 33856
rect 298468 33804 298520 33856
rect 358820 33804 358872 33856
rect 383108 33804 383160 33856
rect 383568 33804 383620 33856
rect 384948 33804 385000 33856
rect 444380 33804 444432 33856
rect 449716 33804 449768 33856
rect 509240 33804 509292 33856
rect 144736 33736 144788 33788
rect 205640 33736 205692 33788
rect 270408 33736 270460 33788
rect 331220 33736 331272 33788
rect 338028 33736 338080 33788
rect 398932 33736 398984 33788
rect 502156 33736 502208 33788
rect 563152 33736 563204 33788
rect 266544 32512 266596 32564
rect 327080 32512 327132 32564
rect 142068 32444 142120 32496
rect 201500 32444 201552 32496
rect 202788 32444 202840 32496
rect 262220 32444 262272 32496
rect 295248 32444 295300 32496
rect 356152 32444 356204 32496
rect 373908 32444 373960 32496
rect 433340 32444 433392 32496
rect 445668 32444 445720 32496
rect 505100 32444 505152 32496
rect 110328 32376 110380 32428
rect 169760 32376 169812 32428
rect 170956 32376 171008 32428
rect 230480 32376 230532 32428
rect 234528 32376 234580 32428
rect 295340 32376 295392 32428
rect 327264 32376 327316 32428
rect 387800 32376 387852 32428
rect 420828 32376 420880 32428
rect 480260 32376 480312 32428
rect 495348 32376 495400 32428
rect 554872 32376 554924 32428
rect 135168 31152 135220 31204
rect 194600 31152 194652 31204
rect 106188 31084 106240 31136
rect 167092 31084 167144 31136
rect 198648 31084 198700 31136
rect 259460 31084 259512 31136
rect 263508 31084 263560 31136
rect 322940 31084 322992 31136
rect 324228 31084 324280 31136
rect 383660 31084 383712 31136
rect 492588 31084 492640 31136
rect 552020 31084 552072 31136
rect 166908 31016 166960 31068
rect 227812 31016 227864 31068
rect 231676 31016 231728 31068
rect 291200 31016 291252 31068
rect 292488 31016 292540 31068
rect 351920 31016 351972 31068
rect 371056 31016 371108 31068
rect 430580 31016 430632 31068
rect 441436 31016 441488 31068
rect 502432 31016 502484 31068
rect 523868 30268 523920 30320
rect 580172 30268 580224 30320
rect 191748 29792 191800 29844
rect 252652 29792 252704 29844
rect 131028 29724 131080 29776
rect 191840 29724 191892 29776
rect 256608 29724 256660 29776
rect 316040 29724 316092 29776
rect 102048 29656 102100 29708
rect 162860 29656 162912 29708
rect 223396 29656 223448 29708
rect 284300 29656 284352 29708
rect 406936 29656 406988 29708
rect 466460 29656 466512 29708
rect 162676 29588 162728 29640
rect 223580 29588 223632 29640
rect 284116 29588 284168 29640
rect 345020 29588 345072 29640
rect 354496 29588 354548 29640
rect 415400 29588 415452 29640
rect 438768 29588 438820 29640
rect 498200 29588 498252 29640
rect 434812 29019 434864 29028
rect 434812 28985 434821 29019
rect 434821 28985 434855 29019
rect 434855 28985 434864 29019
rect 434812 28976 434864 28985
rect 383292 28908 383344 28960
rect 272524 28296 272576 28348
rect 331312 28296 331364 28348
rect 378048 28296 378100 28348
rect 437480 28296 437532 28348
rect 488448 28296 488500 28348
rect 547880 28296 547932 28348
rect 97908 28228 97960 28280
rect 158812 28228 158864 28280
rect 165528 28228 165580 28280
rect 226340 28228 226392 28280
rect 244188 28228 244240 28280
rect 305092 28228 305144 28280
rect 329748 28228 329800 28280
rect 390560 28228 390612 28280
rect 434628 28228 434680 28280
rect 494152 28228 494204 28280
rect 398840 27548 398892 27600
rect 398932 27548 398984 27600
rect 275836 26936 275888 26988
rect 335360 26936 335412 26988
rect 353208 26936 353260 26988
rect 431868 26936 431920 26988
rect 491300 26936 491352 26988
rect 93768 26868 93820 26920
rect 154580 26868 154632 26920
rect 158628 26868 158680 26920
rect 218152 26868 218204 26920
rect 237288 26868 237340 26920
rect 296812 26868 296864 26920
rect 311808 26868 311860 26920
rect 372712 26868 372764 26920
rect 409788 26868 409840 26920
rect 469220 26868 469272 26920
rect 485596 26868 485648 26920
rect 545120 26868 545172 26920
rect 317328 25576 317380 25628
rect 376760 25576 376812 25628
rect 427728 25576 427780 25628
rect 487160 25576 487212 25628
rect 91008 25508 91060 25560
rect 150532 25508 150584 25560
rect 154488 25508 154540 25560
rect 215300 25508 215352 25560
rect 226248 25508 226300 25560
rect 287152 25508 287204 25560
rect 293776 25508 293828 25560
rect 354680 25508 354732 25560
rect 362776 25508 362828 25560
rect 423680 25508 423732 25560
rect 477408 25508 477460 25560
rect 536840 25508 536892 25560
rect 285588 24148 285640 24200
rect 346400 24148 346452 24200
rect 474648 24148 474700 24200
rect 534080 24148 534132 24200
rect 86868 24080 86920 24132
rect 147680 24080 147732 24132
rect 151728 24080 151780 24132
rect 211160 24080 211212 24132
rect 212448 24080 212500 24132
rect 271880 24080 271932 24132
rect 275928 24080 275980 24132
rect 336740 24080 336792 24132
rect 344836 24080 344888 24132
rect 404360 24080 404412 24132
rect 423496 24080 423548 24132
rect 484400 24080 484452 24132
rect 278688 22788 278740 22840
rect 339500 22788 339552 22840
rect 467748 22788 467800 22840
rect 527180 22788 527232 22840
rect 84016 22720 84068 22772
rect 143540 22720 143592 22772
rect 147588 22720 147640 22772
rect 208400 22720 208452 22772
rect 215116 22720 215168 22772
rect 276020 22720 276072 22772
rect 286968 22720 287020 22772
rect 347872 22720 347924 22772
rect 351828 22720 351880 22772
rect 411260 22720 411312 22772
rect 412548 22720 412600 22772
rect 471980 22720 472032 22772
rect 383476 22015 383528 22024
rect 383476 21981 383485 22015
rect 383485 21981 383519 22015
rect 383519 21981 383528 22015
rect 383476 21972 383528 21981
rect 419448 21428 419500 21480
rect 478880 21428 478932 21480
rect 79968 21360 80020 21412
rect 140780 21360 140832 21412
rect 144828 21360 144880 21412
rect 204260 21360 204312 21412
rect 205548 21360 205600 21412
rect 264980 21360 265032 21412
rect 269028 21360 269080 21412
rect 329840 21360 329892 21412
rect 336556 21360 336608 21412
rect 397460 21360 397512 21412
rect 470508 21360 470560 21412
rect 529940 21360 529992 21412
rect 456708 20000 456760 20052
rect 516140 20000 516192 20052
rect 75828 19932 75880 19984
rect 136640 19932 136692 19984
rect 140688 19932 140740 19984
rect 201592 19932 201644 19984
rect 208308 19932 208360 19984
rect 269120 19932 269172 19984
rect 273168 19932 273220 19984
rect 332600 19932 332652 19984
rect 333888 19932 333940 19984
rect 393320 19932 393372 19984
rect 405648 19932 405700 19984
rect 465080 19932 465132 19984
rect 506388 19932 506440 19984
rect 565820 19932 565872 19984
rect 412640 19363 412692 19372
rect 412640 19329 412649 19363
rect 412649 19329 412683 19363
rect 412683 19329 412692 19363
rect 412640 19320 412692 19329
rect 372620 19295 372672 19304
rect 372620 19261 372629 19295
rect 372629 19261 372663 19295
rect 372663 19261 372672 19295
rect 372620 19252 372672 19261
rect 390376 19252 390428 19304
rect 390560 19252 390612 19304
rect 434812 19295 434864 19304
rect 434812 19261 434821 19295
rect 434821 19261 434855 19295
rect 434855 19261 434864 19295
rect 434812 19252 434864 19261
rect 467104 18640 467156 18692
rect 520372 18640 520424 18692
rect 73068 18572 73120 18624
rect 132592 18572 132644 18624
rect 136456 18572 136508 18624
rect 197360 18572 197412 18624
rect 201408 18572 201460 18624
rect 262312 18572 262364 18624
rect 266268 18572 266320 18624
rect 325700 18572 325752 18624
rect 326988 18572 327040 18624
rect 386420 18572 386472 18624
rect 408408 18572 408460 18624
rect 467840 18572 467892 18624
rect 510528 18572 510580 18624
rect 569960 18572 570012 18624
rect 523776 17892 523828 17944
rect 580080 17892 580132 17944
rect 70308 17280 70360 17332
rect 131120 17280 131172 17332
rect 401508 17280 401560 17332
rect 460940 17280 460992 17332
rect 129648 17212 129700 17264
rect 190460 17212 190512 17264
rect 197176 17212 197228 17264
rect 258080 17212 258132 17264
rect 262128 17212 262180 17264
rect 321652 17212 321704 17264
rect 322848 17212 322900 17264
rect 382372 17212 382424 17264
rect 452568 17212 452620 17264
rect 512092 17212 512144 17264
rect 126796 15920 126848 15972
rect 186320 15920 186372 15972
rect 315948 15920 316000 15972
rect 375380 15920 375432 15972
rect 424968 15920 425020 15972
rect 485780 15920 485832 15972
rect 66904 15852 66956 15904
rect 126980 15852 127032 15904
rect 194508 15852 194560 15904
rect 253940 15852 253992 15904
rect 257896 15852 257948 15904
rect 318800 15852 318852 15904
rect 397368 15852 397420 15904
rect 458180 15852 458232 15904
rect 469128 15852 469180 15904
rect 528652 15852 528704 15904
rect 81348 14492 81400 14544
rect 140872 14492 140924 14544
rect 309048 14492 309100 14544
rect 368480 14492 368532 14544
rect 395988 14492 396040 14544
rect 455420 14492 455472 14544
rect 122748 14424 122800 14476
rect 183652 14424 183704 14476
rect 187608 14424 187660 14476
rect 247040 14424 247092 14476
rect 251088 14424 251140 14476
rect 311900 14424 311952 14476
rect 344928 14424 344980 14476
rect 405740 14424 405792 14476
rect 448428 14424 448480 14476
rect 507860 14424 507912 14476
rect 509148 14424 509200 14476
rect 568580 14424 568632 14476
rect 84108 13132 84160 13184
rect 144920 13132 144972 13184
rect 248328 13132 248380 13184
rect 307760 13132 307812 13184
rect 367744 13132 367796 13184
rect 394700 13132 394752 13184
rect 444288 13132 444340 13184
rect 503720 13132 503772 13184
rect 118516 13064 118568 13116
rect 179420 13064 179472 13116
rect 183468 13064 183520 13116
rect 244372 13064 244424 13116
rect 304908 13064 304960 13116
rect 365812 13064 365864 13116
rect 389088 13064 389140 13116
rect 448520 13064 448572 13116
rect 505008 13064 505060 13116
rect 564440 13064 564492 13116
rect 383292 12384 383344 12436
rect 383476 12384 383528 12436
rect 401600 12384 401652 12436
rect 402520 12384 402572 12436
rect 404360 12384 404412 12436
rect 404912 12384 404964 12436
rect 372804 12248 372856 12300
rect 331128 11772 331180 11824
rect 391848 11772 391900 11824
rect 441528 11772 441580 11824
rect 500960 11772 501012 11824
rect 115848 11704 115900 11756
rect 175372 11704 175424 11756
rect 179236 11704 179288 11756
rect 240140 11704 240192 11756
rect 241428 11704 241480 11756
rect 300860 11704 300912 11756
rect 302148 11704 302200 11756
rect 361580 11704 361632 11756
rect 380716 11704 380768 11756
rect 441620 11704 441672 11756
rect 499488 11704 499540 11756
rect 558920 11704 558972 11756
rect 311164 10412 311216 10464
rect 370412 10412 370464 10464
rect 176568 10344 176620 10396
rect 236092 10344 236144 10396
rect 298008 10344 298060 10396
rect 357440 10344 357492 10396
rect 416688 10344 416740 10396
rect 477592 10344 477644 10396
rect 111708 10276 111760 10328
rect 172520 10276 172572 10328
rect 233148 10276 233200 10328
rect 293960 10276 294012 10328
rect 355968 10276 356020 10328
rect 416872 10276 416924 10328
rect 437388 10276 437440 10328
rect 496820 10276 496872 10328
rect 498108 10276 498160 10328
rect 557540 10276 557592 10328
rect 434812 9775 434864 9784
rect 434812 9741 434821 9775
rect 434821 9741 434855 9775
rect 434855 9741 434864 9775
rect 434812 9732 434864 9741
rect 390652 9596 390704 9648
rect 411260 9596 411312 9648
rect 415400 9596 415452 9648
rect 434812 9596 434864 9648
rect 390652 9460 390704 9512
rect 230388 8984 230440 9036
rect 290740 8984 290792 9036
rect 291108 8984 291160 9036
rect 351368 8984 351420 9036
rect 108948 8916 109000 8968
rect 169392 8916 169444 8968
rect 172428 8916 172480 8968
rect 233700 8916 233752 8968
rect 347688 8916 347740 8968
rect 408592 8916 408644 8968
rect 430488 8916 430540 8968
rect 490564 8916 490616 8968
rect 491208 8916 491260 8968
rect 551192 8916 551244 8968
rect 137928 7624 137980 7676
rect 199200 7624 199252 7676
rect 223488 7624 223540 7676
rect 283656 7624 283708 7676
rect 340788 7624 340840 7676
rect 401324 7624 401376 7676
rect 433340 7624 433392 7676
rect 434628 7624 434680 7676
rect 481548 7624 481600 7676
rect 541716 7624 541768 7676
rect 104808 7556 104860 7608
rect 165896 7556 165948 7608
rect 169668 7556 169720 7608
rect 230112 7556 230164 7608
rect 284208 7556 284260 7608
rect 344284 7556 344336 7608
rect 382372 7556 382424 7608
rect 383568 7556 383620 7608
rect 408500 7556 408552 7608
rect 409696 7556 409748 7608
rect 426348 7556 426400 7608
rect 486976 7556 487028 7608
rect 162768 6264 162820 6316
rect 222936 6264 222988 6316
rect 219348 6196 219400 6248
rect 279976 6196 280028 6248
rect 282828 6196 282880 6248
rect 343088 6196 343140 6248
rect 423588 6196 423640 6248
rect 483480 6196 483532 6248
rect 100576 6128 100628 6180
rect 162308 6128 162360 6180
rect 209688 6128 209740 6180
rect 270592 6128 270644 6180
rect 280068 6128 280120 6180
rect 340696 6128 340748 6180
rect 345664 6128 345716 6180
rect 379980 6128 380032 6180
rect 398748 6128 398800 6180
rect 459652 6128 459704 6180
rect 516048 6128 516100 6180
rect 576216 6128 576268 6180
rect 380808 5448 380860 5500
rect 440608 5448 440660 5500
rect 369768 5380 369820 5432
rect 429936 5380 429988 5432
rect 455328 5380 455380 5432
rect 515588 5380 515640 5432
rect 365628 5312 365680 5364
rect 426348 5312 426400 5364
rect 459468 5312 459520 5364
rect 519084 5312 519136 5364
rect 387708 5244 387760 5296
rect 447784 5244 447836 5296
rect 462228 5244 462280 5296
rect 522672 5244 522724 5296
rect 376668 5176 376720 5228
rect 437020 5176 437072 5228
rect 466368 5176 466420 5228
rect 526260 5176 526312 5228
rect 358728 5108 358780 5160
rect 419172 5108 419224 5160
rect 473268 5108 473320 5160
rect 533436 5108 533488 5160
rect 394608 5040 394660 5092
rect 454868 5040 454920 5092
rect 480168 5040 480220 5092
rect 540520 5040 540572 5092
rect 362868 4972 362920 5024
rect 422760 4972 422812 5024
rect 484308 4972 484360 5024
rect 544108 4972 544160 5024
rect 133788 4904 133840 4956
rect 194416 4904 194468 4956
rect 255228 4904 255280 4956
rect 315764 4904 315816 4956
rect 383292 4904 383344 4956
rect 444196 4904 444248 4956
rect 463608 4904 463660 4956
rect 523868 4904 523920 4956
rect 66168 4836 66220 4888
rect 126612 4836 126664 4888
rect 190368 4836 190420 4888
rect 251456 4836 251508 4888
rect 303528 4836 303580 4888
rect 364524 4836 364576 4888
rect 390468 4836 390520 4888
rect 68928 4768 68980 4820
rect 130200 4768 130252 4820
rect 173808 4768 173860 4820
rect 234804 4768 234856 4820
rect 252468 4768 252520 4820
rect 313372 4768 313424 4820
rect 372528 4768 372580 4820
rect 425060 4768 425112 4820
rect 487068 4836 487120 4888
rect 547696 4836 547748 4888
rect 476028 4768 476080 4820
rect 536932 4768 536984 4820
rect 451372 4700 451424 4752
rect 528652 4156 528704 4208
rect 529848 4156 529900 4208
rect 118608 4088 118660 4140
rect 178960 4088 179012 4140
rect 179328 4088 179380 4140
rect 239588 4088 239640 4140
rect 264888 4088 264940 4140
rect 325240 4088 325292 4140
rect 379428 4088 379480 4140
rect 439412 4088 439464 4140
rect 442908 4088 442960 4140
rect 503628 4088 503680 4140
rect 514668 4088 514720 4140
rect 575020 4088 575072 4140
rect 150348 4020 150400 4072
rect 211068 4020 211120 4072
rect 240048 4020 240100 4072
rect 300308 4020 300360 4072
rect 350448 4020 350500 4072
rect 410892 4020 410944 4072
rect 411168 4020 411220 4072
rect 471520 4020 471572 4072
rect 493968 4020 494020 4072
rect 553584 4020 553636 4072
rect 143448 3952 143500 4004
rect 203892 3952 203944 4004
rect 231768 3952 231820 4004
rect 246948 3952 247000 4004
rect 307392 3952 307444 4004
rect 318708 3952 318760 4004
rect 378784 3952 378836 4004
rect 386328 3952 386380 4004
rect 446588 3952 446640 4004
rect 496728 3952 496780 4004
rect 557172 3952 557224 4004
rect 88248 3884 88300 3936
rect 149244 3884 149296 3936
rect 161388 3884 161440 3936
rect 221740 3884 221792 3936
rect 229008 3884 229060 3936
rect 289544 3884 289596 3936
rect 300768 3884 300820 3936
rect 360936 3884 360988 3936
rect 393228 3884 393280 3936
rect 453672 3884 453724 3936
rect 500868 3884 500920 3936
rect 560760 3884 560812 3936
rect 128268 3816 128320 3868
rect 189632 3816 189684 3868
rect 197268 3816 197320 3868
rect 257436 3816 257488 3868
rect 257988 3816 258040 3868
rect 318064 3816 318116 3868
rect 325608 3816 325660 3868
rect 385868 3816 385920 3868
rect 400128 3816 400180 3868
rect 460756 3816 460808 3868
rect 503444 3816 503496 3868
rect 564348 3816 564400 3868
rect 114468 3748 114520 3800
rect 175280 3748 175332 3800
rect 200028 3748 200080 3800
rect 261024 3748 261076 3800
rect 262220 3748 262272 3800
rect 263416 3748 263468 3800
rect 289728 3748 289780 3800
rect 350264 3748 350316 3800
rect 354588 3748 354640 3800
rect 414480 3748 414532 3800
rect 447048 3748 447100 3800
rect 507216 3748 507268 3800
rect 513288 3748 513340 3800
rect 573824 3748 573876 3800
rect 121368 3680 121420 3732
rect 182548 3680 182600 3732
rect 201500 3680 201552 3732
rect 202696 3680 202748 3732
rect 206928 3680 206980 3732
rect 268108 3680 268160 3732
rect 296628 3680 296680 3732
rect 357348 3680 357400 3732
rect 361488 3680 361540 3732
rect 421564 3680 421616 3732
rect 422208 3680 422260 3732
rect 482284 3680 482336 3732
rect 511908 3680 511960 3732
rect 571340 3680 571392 3732
rect 71688 3612 71740 3664
rect 132500 3612 132552 3664
rect 153108 3612 153160 3664
rect 214656 3612 214708 3664
rect 235908 3612 235960 3664
rect 296720 3612 296772 3664
rect 321652 3612 321704 3664
rect 322848 3612 322900 3664
rect 328368 3612 328420 3664
rect 389456 3612 389508 3664
rect 418068 3612 418120 3664
rect 478696 3612 478748 3664
rect 507768 3612 507820 3664
rect 567844 3612 567896 3664
rect 78588 3544 78640 3596
rect 139676 3544 139728 3596
rect 140872 3544 140924 3596
rect 142068 3544 142120 3596
rect 150532 3544 150584 3596
rect 151544 3544 151596 3596
rect 157248 3544 157300 3596
rect 218060 3544 218112 3596
rect 218152 3544 218204 3596
rect 219348 3544 219400 3596
rect 236092 3544 236144 3596
rect 237196 3544 237248 3596
rect 293132 3544 293184 3596
rect 305000 3544 305052 3596
rect 306196 3544 306248 3596
rect 310428 3544 310480 3596
rect 368020 3544 368072 3596
rect 415308 3544 415360 3596
rect 475108 3544 475160 3596
rect 494152 3544 494204 3596
rect 495348 3544 495400 3596
rect 517428 3544 517480 3596
rect 577412 3544 577464 3596
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 74356 3476 74408 3528
rect 132592 3476 132644 3528
rect 133788 3476 133840 3528
rect 171048 3476 171100 3528
rect 232504 3476 232556 3528
rect 244280 3476 244332 3528
rect 245568 3476 245620 3528
rect 249708 3476 249760 3528
rect 310980 3476 311032 3528
rect 321468 3476 321520 3528
rect 382372 3476 382424 3528
rect 429108 3476 429160 3528
rect 489368 3476 489420 3528
rect 518808 3476 518860 3528
rect 578608 3476 578660 3528
rect 572 3408 624 3460
rect 62120 3408 62172 3460
rect 95148 3408 95200 3460
rect 156328 3408 156380 3460
rect 164148 3408 164200 3460
rect 225328 3408 225380 3460
rect 242808 3408 242860 3460
rect 303804 3408 303856 3460
rect 307668 3408 307720 3460
rect 365720 3408 365772 3460
rect 366916 3408 366968 3460
rect 371148 3408 371200 3460
rect 432328 3408 432380 3460
rect 436008 3408 436060 3460
rect 496544 3408 496596 3460
rect 521568 3408 521620 3460
rect 582196 3408 582248 3460
rect 125508 3340 125560 3392
rect 183560 3340 183612 3392
rect 184848 3340 184900 3392
rect 204168 3340 204220 3392
rect 264612 3340 264664 3392
rect 270500 3340 270552 3392
rect 271696 3340 271748 3392
rect 287060 3340 287112 3392
rect 288348 3340 288400 3392
rect 293868 3340 293920 3392
rect 353760 3340 353812 3392
rect 357164 3340 357216 3392
rect 417976 3340 418028 3392
rect 451280 3340 451332 3392
rect 452476 3340 452528 3392
rect 467840 3340 467892 3392
rect 469128 3340 469180 3392
rect 471888 3340 471940 3392
rect 532240 3340 532292 3392
rect 536840 3340 536892 3392
rect 538128 3340 538180 3392
rect 571432 3340 571484 3392
rect 572628 3340 572680 3392
rect 136088 3272 136140 3324
rect 136548 3272 136600 3324
rect 196808 3272 196860 3324
rect 215208 3272 215260 3324
rect 275284 3272 275336 3324
rect 343548 3272 343600 3324
rect 403716 3272 403768 3324
rect 478788 3272 478840 3324
rect 539324 3272 539376 3324
rect 100668 3204 100720 3256
rect 161112 3204 161164 3256
rect 175372 3204 175424 3256
rect 176568 3204 176620 3256
rect 186044 3204 186096 3256
rect 193128 3204 193180 3256
rect 253848 3204 253900 3256
rect 314660 3204 314712 3256
rect 375196 3204 375248 3256
rect 460848 3204 460900 3256
rect 521476 3204 521528 3256
rect 107568 3136 107620 3188
rect 168196 3136 168248 3188
rect 186228 3136 186280 3188
rect 246764 3136 246816 3188
rect 332508 3136 332560 3188
rect 393044 3136 393096 3188
rect 453948 3136 454000 3188
rect 514392 3136 514444 3188
rect 92388 3068 92440 3120
rect 152740 3068 152792 3120
rect 222108 3068 222160 3120
rect 282460 3068 282512 3120
rect 336648 3068 336700 3120
rect 396632 3068 396684 3120
rect 458088 3068 458140 3120
rect 517888 3068 517940 3120
rect 99288 3000 99340 3052
rect 159916 3000 159968 3052
rect 371608 3000 371660 3052
rect 464988 3000 465040 3052
rect 525064 3000 525116 3052
rect 440148 2932 440200 2984
rect 500132 2932 500184 2984
rect 433156 2864 433208 2916
rect 492956 2864 493008 2916
rect 393320 2796 393372 2848
rect 394700 2796 394752 2848
rect 397460 2796 397512 2848
rect 412640 2796 412692 2848
rect 419540 2796 419592 2848
rect 426440 2796 426492 2848
rect 427912 2796 427964 2848
rect 430580 2796 430632 2848
rect 394240 2728 394292 2780
rect 395436 2728 395488 2780
rect 397828 2728 397880 2780
rect 413284 2728 413336 2780
rect 420368 2728 420420 2780
rect 427544 2728 427596 2780
rect 428740 2728 428792 2780
rect 431132 2728 431184 2780
rect 347780 2048 347832 2100
rect 349068 2048 349120 2100
rect 375380 552 375432 604
rect 376392 552 376444 604
rect 376760 552 376812 604
rect 377588 552 377640 604
rect 383660 552 383712 604
rect 384672 552 384724 604
rect 386420 552 386472 604
rect 387064 552 387116 604
rect 387800 552 387852 604
rect 388260 552 388312 604
rect 405740 552 405792 604
rect 406108 552 406160 604
rect 412088 595 412140 604
rect 412088 561 412097 595
rect 412097 561 412131 595
rect 412131 561 412140 595
rect 412088 552 412140 561
rect 415676 595 415728 604
rect 415676 561 415685 595
rect 415685 561 415719 595
rect 415719 561 415728 595
rect 415676 552 415728 561
rect 435824 595 435876 604
rect 435824 561 435833 595
rect 435833 561 435867 595
rect 435867 561 435876 595
rect 435824 552 435876 561
rect 455420 552 455472 604
rect 456064 552 456116 604
rect 456892 552 456944 604
rect 457260 552 457312 604
rect 471980 552 472032 604
rect 472716 552 472768 604
rect 473360 552 473412 604
rect 473912 552 473964 604
rect 478880 552 478932 604
rect 479892 552 479944 604
rect 579620 552 579672 604
rect 579804 552 579856 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703474 73016 703520
rect 72804 703446 73016 703474
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3422 682272 3478 682281
rect 3422 682207 3478 682216
rect 3436 636206 3464 682207
rect 8128 679046 8156 685850
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 3514 667992 3570 668001
rect 3514 667927 3570 667936
rect 3424 636200 3476 636206
rect 3424 636142 3476 636148
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 593366 3464 624815
rect 3528 622402 3556 667927
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654158 8064 663734
rect 8024 654152 8076 654158
rect 8024 654094 8076 654100
rect 8208 654152 8260 654158
rect 8208 654094 8260 654100
rect 3606 653576 3662 653585
rect 3606 653511 3662 653520
rect 3516 622396 3568 622402
rect 3516 622338 3568 622344
rect 3514 610464 3570 610473
rect 3514 610399 3570 610408
rect 3424 593360 3476 593366
rect 3424 593302 3476 593308
rect 3528 579630 3556 610399
rect 3620 608598 3648 653511
rect 8220 645318 8248 654094
rect 8208 645312 8260 645318
rect 8208 645254 8260 645260
rect 24780 645182 24808 699654
rect 41340 645250 41368 700334
rect 72804 698306 72832 703446
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 703474 137876 703520
rect 137756 703446 137876 703474
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 72712 698278 72832 698306
rect 72712 694142 72740 698278
rect 72700 694136 72752 694142
rect 72700 694078 72752 694084
rect 72516 684616 72568 684622
rect 72516 684558 72568 684564
rect 72528 684486 72556 684558
rect 72516 684480 72568 684486
rect 72516 684422 72568 684428
rect 72792 676116 72844 676122
rect 72792 676058 72844 676064
rect 72804 669390 72832 676058
rect 72792 669384 72844 669390
rect 72792 669326 72844 669332
rect 72792 669248 72844 669254
rect 72792 669190 72844 669196
rect 72804 659682 72832 669190
rect 72804 659654 73016 659682
rect 72988 650026 73016 659654
rect 72988 649998 73108 650026
rect 73080 645386 73108 649998
rect 73068 645380 73120 645386
rect 73068 645322 73120 645328
rect 89640 645318 89668 699654
rect 70492 645312 70544 645318
rect 70492 645254 70544 645260
rect 89628 645312 89680 645318
rect 89628 645254 89680 645260
rect 41328 645244 41380 645250
rect 41328 645186 41380 645192
rect 24768 645176 24820 645182
rect 24768 645118 24820 645124
rect 70504 643076 70532 645254
rect 104532 645244 104584 645250
rect 104532 645186 104584 645192
rect 87512 645176 87564 645182
rect 87512 645118 87564 645124
rect 87524 643076 87552 645118
rect 104544 643076 104572 645186
rect 106200 645182 106228 699654
rect 137756 698290 137784 703446
rect 137744 698284 137796 698290
rect 137744 698226 137796 698232
rect 137928 698284 137980 698290
rect 137928 698226 137980 698232
rect 137940 695502 137968 698226
rect 154132 695570 154160 703520
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 137928 695496 137980 695502
rect 137928 695438 137980 695444
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 137836 685908 137888 685914
rect 137836 685850 137888 685856
rect 137848 679046 137876 685850
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 137836 679040 137888 679046
rect 137836 678982 137888 678988
rect 137744 678972 137796 678978
rect 137744 678914 137796 678920
rect 137756 673538 137784 678914
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 137744 673532 137796 673538
rect 137744 673474 137796 673480
rect 137928 673532 137980 673538
rect 137928 673474 137980 673480
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 137940 663762 137968 673474
rect 154500 663762 154528 673474
rect 137756 663734 137968 663762
rect 154316 663734 154528 663762
rect 137756 654158 137784 663734
rect 154316 654158 154344 663734
rect 137744 654152 137796 654158
rect 137744 654094 137796 654100
rect 137928 654152 137980 654158
rect 137928 654094 137980 654100
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 137940 645386 137968 654094
rect 121552 645380 121604 645386
rect 121552 645322 121604 645328
rect 137928 645380 137980 645386
rect 137928 645322 137980 645328
rect 106188 645176 106240 645182
rect 106188 645118 106240 645124
rect 121564 643076 121592 645322
rect 138572 645312 138624 645318
rect 138572 645254 138624 645260
rect 138584 643076 138612 645254
rect 154500 645250 154528 654094
rect 154488 645244 154540 645250
rect 154488 645186 154540 645192
rect 171060 645182 171088 700198
rect 172704 645380 172756 645386
rect 172704 645322 172756 645328
rect 155592 645176 155644 645182
rect 155592 645118 155644 645124
rect 171048 645176 171100 645182
rect 171048 645118 171100 645124
rect 155604 643076 155632 645118
rect 172716 643076 172744 645322
rect 202800 645250 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 678994 219112 685850
rect 218992 678966 219112 678994
rect 218992 676190 219020 678966
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 219084 659682 219112 666538
rect 219084 659654 219296 659682
rect 219268 650026 219296 659654
rect 219268 649998 219388 650026
rect 189724 645244 189776 645250
rect 189724 645186 189776 645192
rect 202788 645244 202840 645250
rect 202788 645186 202840 645192
rect 189736 643076 189764 645186
rect 219360 645182 219388 649998
rect 235920 645250 235948 699654
rect 223764 645244 223816 645250
rect 223764 645186 223816 645192
rect 235908 645244 235960 645250
rect 235908 645186 235960 645192
rect 257896 645244 257948 645250
rect 257896 645186 257948 645192
rect 206744 645176 206796 645182
rect 206744 645118 206796 645124
rect 219348 645176 219400 645182
rect 219348 645118 219400 645124
rect 206756 643076 206784 645118
rect 223776 643076 223804 645186
rect 240784 645176 240836 645182
rect 240784 645118 240836 645124
rect 240796 643076 240824 645118
rect 257908 643076 257936 645186
rect 267660 645182 267688 703520
rect 283852 695570 283880 703520
rect 300136 699718 300164 703520
rect 332520 699718 332548 703520
rect 348804 700330 348832 703520
rect 344284 700324 344336 700330
rect 344284 700266 344336 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 326988 699712 327040 699718
rect 326988 699654 327040 699660
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 283840 695564 283892 695570
rect 283840 695506 283892 695512
rect 283932 695564 283984 695570
rect 283932 695506 283984 695512
rect 283944 688634 283972 695506
rect 283932 688628 283984 688634
rect 283932 688570 283984 688576
rect 284116 688628 284168 688634
rect 284116 688570 284168 688576
rect 284128 685846 284156 688570
rect 284116 685840 284168 685846
rect 284116 685782 284168 685788
rect 284024 676252 284076 676258
rect 284024 676194 284076 676200
rect 284036 673538 284064 676194
rect 284024 673532 284076 673538
rect 284024 673474 284076 673480
rect 284208 673532 284260 673538
rect 284208 673474 284260 673480
rect 284220 663762 284248 673474
rect 284036 663734 284248 663762
rect 284036 654158 284064 663734
rect 284024 654152 284076 654158
rect 284024 654094 284076 654100
rect 284208 654152 284260 654158
rect 284208 654094 284260 654100
rect 284220 645182 284248 654094
rect 267648 645176 267700 645182
rect 267648 645118 267700 645124
rect 274916 645176 274968 645182
rect 274916 645118 274968 645124
rect 284208 645176 284260 645182
rect 284208 645118 284260 645124
rect 291936 645176 291988 645182
rect 291936 645118 291988 645124
rect 274928 643076 274956 645118
rect 291948 643076 291976 645118
rect 300780 644910 300808 699654
rect 327000 645522 327028 699654
rect 344296 645862 344324 700266
rect 364996 699718 365024 703520
rect 394608 700460 394660 700466
rect 394608 700402 394660 700408
rect 378048 700324 378100 700330
rect 378048 700266 378100 700272
rect 360108 699712 360160 699718
rect 360108 699654 360160 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 342996 645856 343048 645862
rect 342996 645798 343048 645804
rect 344284 645856 344336 645862
rect 344284 645798 344336 645804
rect 325976 645516 326028 645522
rect 325976 645458 326028 645464
rect 326988 645516 327040 645522
rect 326988 645458 327040 645464
rect 300768 644904 300820 644910
rect 300768 644846 300820 644852
rect 308956 644904 309008 644910
rect 308956 644846 309008 644852
rect 308968 643076 308996 644846
rect 325988 643076 326016 645458
rect 343008 643076 343036 645798
rect 360120 643076 360148 699654
rect 378060 645862 378088 700266
rect 377128 645856 377180 645862
rect 377128 645798 377180 645804
rect 378048 645856 378100 645862
rect 378048 645798 378100 645804
rect 377140 643076 377168 645798
rect 394620 642954 394648 700402
rect 397472 700330 397500 703520
rect 413664 700466 413692 703520
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 429856 700398 429884 703520
rect 411168 700392 411220 700398
rect 411168 700334 411220 700340
rect 429844 700392 429896 700398
rect 429844 700334 429896 700340
rect 445668 700392 445720 700398
rect 445668 700334 445720 700340
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 411180 643076 411208 700334
rect 429108 700324 429160 700330
rect 429108 700266 429160 700272
rect 429120 645862 429148 700266
rect 428188 645856 428240 645862
rect 428188 645798 428240 645804
rect 429108 645856 429160 645862
rect 429108 645798 429160 645804
rect 428200 643076 428228 645798
rect 445680 643090 445708 700334
rect 462332 700330 462360 703520
rect 463608 700460 463660 700466
rect 463608 700402 463660 700408
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 463620 645862 463648 700402
rect 478524 700398 478552 703520
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 514668 700460 514720 700466
rect 514668 700402 514720 700408
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 496728 700392 496780 700398
rect 496728 700334 496780 700340
rect 480168 700324 480220 700330
rect 480168 700266 480220 700272
rect 480180 645862 480208 700266
rect 462320 645856 462372 645862
rect 462320 645798 462372 645804
rect 463608 645856 463660 645862
rect 463608 645798 463660 645804
rect 479340 645856 479392 645862
rect 479340 645798 479392 645804
rect 480168 645856 480220 645862
rect 480168 645798 480220 645804
rect 445326 643062 445708 643090
rect 462332 643076 462360 645798
rect 479352 643076 479380 645798
rect 496740 643090 496768 700334
rect 514680 645658 514708 700402
rect 527192 700330 527220 703520
rect 543476 700398 543504 703520
rect 559668 700466 559696 703520
rect 559656 700460 559708 700466
rect 559656 700402 559708 700408
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 523776 696992 523828 696998
rect 523776 696934 523828 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 523684 685908 523736 685914
rect 523684 685850 523736 685856
rect 513380 645652 513432 645658
rect 513380 645594 513432 645600
rect 514668 645652 514720 645658
rect 514668 645594 514720 645600
rect 496386 643062 496768 643090
rect 513392 643076 513420 645594
rect 394174 642926 394648 642954
rect 59360 636200 59412 636206
rect 59360 636142 59412 636148
rect 59372 636041 59400 636142
rect 59358 636032 59414 636041
rect 59358 635967 59414 635976
rect 523696 623257 523724 685850
rect 523788 636585 523816 696934
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580262 674656 580318 674665
rect 580262 674591 580318 674600
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 523868 638988 523920 638994
rect 523868 638930 523920 638936
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 523774 636576 523830 636585
rect 523774 636511 523830 636520
rect 523682 623248 523738 623257
rect 523682 623183 523738 623192
rect 59360 622396 59412 622402
rect 59360 622338 59412 622344
rect 59372 621761 59400 622338
rect 59358 621752 59414 621761
rect 59358 621687 59414 621696
rect 3608 608592 3660 608598
rect 3608 608534 3660 608540
rect 59360 608592 59412 608598
rect 59360 608534 59412 608540
rect 59372 607481 59400 608534
rect 59358 607472 59414 607481
rect 59358 607407 59414 607416
rect 523776 603152 523828 603158
rect 523776 603094 523828 603100
rect 523684 597508 523736 597514
rect 523684 597450 523736 597456
rect 523696 596601 523724 597450
rect 523682 596592 523738 596601
rect 523682 596527 523738 596536
rect 3606 596048 3662 596057
rect 3606 595983 3662 595992
rect 3516 579624 3568 579630
rect 3516 579566 3568 579572
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 550594 3464 567287
rect 3620 565826 3648 595983
rect 59360 593360 59412 593366
rect 59360 593302 59412 593308
rect 59372 593201 59400 593302
rect 59358 593192 59414 593201
rect 59358 593127 59414 593136
rect 523684 592068 523736 592074
rect 523684 592010 523736 592016
rect 59360 579624 59412 579630
rect 59360 579566 59412 579572
rect 59372 578921 59400 579566
rect 59358 578912 59414 578921
rect 59358 578847 59414 578856
rect 3608 565820 3660 565826
rect 3608 565762 3660 565768
rect 59360 565820 59412 565826
rect 59360 565762 59412 565768
rect 59372 564641 59400 565762
rect 59358 564632 59414 564641
rect 59358 564567 59414 564576
rect 3514 553072 3570 553081
rect 3514 553007 3570 553016
rect 3424 550588 3476 550594
rect 3424 550530 3476 550536
rect 3422 538656 3478 538665
rect 3422 538591 3478 538600
rect 3436 522986 3464 538591
rect 3528 536790 3556 553007
rect 59360 550588 59412 550594
rect 59360 550530 59412 550536
rect 59372 550361 59400 550530
rect 59358 550352 59414 550361
rect 59358 550287 59414 550296
rect 523696 543289 523724 592010
rect 523788 556617 523816 603094
rect 523880 583273 523908 638930
rect 580276 609958 580304 674591
rect 580446 651128 580502 651137
rect 580446 651063 580502 651072
rect 580354 627736 580410 627745
rect 580354 627671 580410 627680
rect 524328 609952 524380 609958
rect 524326 609920 524328 609929
rect 580264 609952 580316 609958
rect 524380 609920 524382 609929
rect 580264 609894 580316 609900
rect 524326 609855 524382 609864
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 523866 583264 523922 583273
rect 523866 583199 523922 583208
rect 580262 580816 580318 580825
rect 580262 580751 580318 580760
rect 524326 569936 524382 569945
rect 524326 569871 524328 569880
rect 524380 569871 524382 569880
rect 524328 569842 524380 569848
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 523774 556608 523830 556617
rect 523774 556543 523830 556552
rect 580184 556238 580212 557223
rect 523868 556232 523920 556238
rect 523868 556174 523920 556180
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 523776 545148 523828 545154
rect 523776 545090 523828 545096
rect 523682 543280 523738 543289
rect 523682 543215 523738 543224
rect 3516 536784 3568 536790
rect 3516 536726 3568 536732
rect 59360 536784 59412 536790
rect 59360 536726 59412 536732
rect 59372 536081 59400 536726
rect 59358 536072 59414 536081
rect 59358 536007 59414 536016
rect 523224 531276 523276 531282
rect 523224 531218 523276 531224
rect 523236 529961 523264 531218
rect 523222 529952 523278 529961
rect 523222 529887 523278 529896
rect 3424 522980 3476 522986
rect 3424 522922 3476 522928
rect 59360 522980 59412 522986
rect 59360 522922 59412 522928
rect 59372 521801 59400 522922
rect 59358 521792 59414 521801
rect 59358 521727 59414 521736
rect 3330 509960 3386 509969
rect 3330 509895 3386 509904
rect 3344 507822 3372 509895
rect 3332 507816 3384 507822
rect 3332 507758 3384 507764
rect 59360 507816 59412 507822
rect 59360 507758 59412 507764
rect 59372 507521 59400 507758
rect 59358 507512 59414 507521
rect 59358 507447 59414 507456
rect 523788 503305 523816 545090
rect 523880 516633 523908 556174
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 580276 531282 580304 580751
rect 580368 569906 580396 627671
rect 580460 597514 580488 651063
rect 580448 597508 580500 597514
rect 580448 597450 580500 597456
rect 580356 569900 580408 569906
rect 580356 569842 580408 569848
rect 580354 533896 580410 533905
rect 580354 533831 580410 533840
rect 580264 531276 580316 531282
rect 580264 531218 580316 531224
rect 523866 516624 523922 516633
rect 523866 516559 523922 516568
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 523868 509312 523920 509318
rect 523868 509254 523920 509260
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 523774 503296 523830 503305
rect 523774 503231 523830 503240
rect 523776 498228 523828 498234
rect 523776 498170 523828 498176
rect 3330 495544 3386 495553
rect 3330 495479 3386 495488
rect 3344 494018 3372 495479
rect 3332 494012 3384 494018
rect 3332 493954 3384 493960
rect 59360 494012 59412 494018
rect 59360 493954 59412 493960
rect 59372 493241 59400 493954
rect 59358 493232 59414 493241
rect 59358 493167 59414 493176
rect 523684 485852 523736 485858
rect 523684 485794 523736 485800
rect 3606 481128 3662 481137
rect 3606 481063 3662 481072
rect 3620 480214 3648 481063
rect 3608 480208 3660 480214
rect 3608 480150 3660 480156
rect 59360 480208 59412 480214
rect 59360 480150 59412 480156
rect 59372 478961 59400 480150
rect 59358 478952 59414 478961
rect 59358 478887 59414 478896
rect 59358 464672 59414 464681
rect 59358 464607 59414 464616
rect 59372 463758 59400 464607
rect 3424 463752 3476 463758
rect 3424 463694 3476 463700
rect 59360 463752 59412 463758
rect 59360 463694 59412 463700
rect 3436 452441 3464 463694
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 59358 450392 59414 450401
rect 59358 450327 59414 450336
rect 59372 449954 59400 450327
rect 523696 449993 523724 485794
rect 523788 463321 523816 498170
rect 523880 476649 523908 509254
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 580368 491298 580396 533831
rect 524328 491292 524380 491298
rect 524328 491234 524380 491240
rect 580356 491292 580408 491298
rect 580356 491234 580408 491240
rect 524340 489977 524368 491234
rect 524326 489968 524382 489977
rect 524326 489903 524382 489912
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 523866 476640 523922 476649
rect 523866 476575 523922 476584
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 523774 463312 523830 463321
rect 523774 463247 523830 463256
rect 580184 462398 580212 463383
rect 523868 462392 523920 462398
rect 523868 462334 523920 462340
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 523776 451308 523828 451314
rect 523776 451250 523828 451256
rect 523682 449984 523738 449993
rect 3424 449948 3476 449954
rect 3424 449890 3476 449896
rect 59360 449948 59412 449954
rect 523682 449919 523738 449928
rect 59360 449890 59412 449896
rect 3436 438025 3464 449890
rect 523684 438932 523736 438938
rect 523684 438874 523736 438880
rect 3422 438016 3478 438025
rect 3422 437951 3478 437960
rect 3424 436144 3476 436150
rect 59360 436144 59412 436150
rect 3424 436086 3476 436092
rect 59358 436112 59360 436121
rect 59412 436112 59414 436121
rect 3436 423745 3464 436086
rect 59358 436047 59414 436056
rect 3422 423736 3478 423745
rect 3422 423671 3478 423680
rect 59358 421832 59414 421841
rect 59358 421767 59414 421776
rect 59372 420986 59400 421767
rect 3516 420980 3568 420986
rect 3516 420922 3568 420928
rect 59360 420980 59412 420986
rect 59360 420922 59412 420928
rect 3424 407176 3476 407182
rect 3424 407118 3476 407124
rect 3436 380633 3464 407118
rect 3528 395049 3556 420922
rect 523696 410009 523724 438874
rect 523788 423337 523816 451250
rect 523880 436665 523908 462334
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580184 451314 580212 451687
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 523866 436656 523922 436665
rect 523866 436591 523922 436600
rect 523774 423328 523830 423337
rect 523774 423263 523830 423272
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 580184 415478 580212 416463
rect 523868 415472 523920 415478
rect 523868 415414 523920 415420
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 523682 410000 523738 410009
rect 523682 409935 523738 409944
rect 59358 407552 59414 407561
rect 59358 407487 59414 407496
rect 59372 407182 59400 407487
rect 59360 407176 59412 407182
rect 59360 407118 59412 407124
rect 523776 404388 523828 404394
rect 523776 404330 523828 404336
rect 3514 395040 3570 395049
rect 3514 394975 3570 394984
rect 59358 393272 59414 393281
rect 59358 393207 59414 393216
rect 59372 392018 59400 393207
rect 3516 392012 3568 392018
rect 3516 391954 3568 391960
rect 59360 392012 59412 392018
rect 59360 391954 59412 391960
rect 523684 392012 523736 392018
rect 523684 391954 523736 391960
rect 3422 380624 3478 380633
rect 3422 380559 3478 380568
rect 3424 378208 3476 378214
rect 3424 378150 3476 378156
rect 3436 337521 3464 378150
rect 3528 366217 3556 391954
rect 59358 378992 59414 379001
rect 59358 378927 59414 378936
rect 59372 378214 59400 378927
rect 59360 378208 59412 378214
rect 59360 378150 59412 378156
rect 523696 370025 523724 391954
rect 523788 383353 523816 404330
rect 523880 396681 523908 415414
rect 580170 404832 580226 404841
rect 580170 404767 580226 404776
rect 580184 404394 580212 404767
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 523866 396672 523922 396681
rect 523866 396607 523922 396616
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 580184 392018 580212 392935
rect 580172 392012 580224 392018
rect 580172 391954 580224 391960
rect 523774 383344 523830 383353
rect 523774 383279 523830 383288
rect 523682 370016 523738 370025
rect 523682 369951 523738 369960
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580184 368558 580212 369543
rect 523684 368552 523736 368558
rect 523684 368494 523736 368500
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 3514 366208 3570 366217
rect 3514 366143 3570 366152
rect 59358 364712 59414 364721
rect 59358 364647 59414 364656
rect 59372 364410 59400 364647
rect 3516 364404 3568 364410
rect 3516 364346 3568 364352
rect 59360 364404 59412 364410
rect 59360 364346 59412 364352
rect 3422 337512 3478 337521
rect 3422 337447 3478 337456
rect 3424 335368 3476 335374
rect 3424 335310 3476 335316
rect 3436 294409 3464 335310
rect 3528 323105 3556 364346
rect 523696 356697 523724 368494
rect 580170 357912 580226 357921
rect 580170 357847 580226 357856
rect 580184 357474 580212 357847
rect 523776 357468 523828 357474
rect 523776 357410 523828 357416
rect 580172 357468 580224 357474
rect 580172 357410 580224 357416
rect 523682 356688 523738 356697
rect 523682 356623 523738 356632
rect 59358 350432 59414 350441
rect 59358 350367 59414 350376
rect 59372 349178 59400 350367
rect 3608 349172 3660 349178
rect 3608 349114 3660 349120
rect 59360 349172 59412 349178
rect 59360 349114 59412 349120
rect 3514 323096 3570 323105
rect 3514 323031 3570 323040
rect 3516 321632 3568 321638
rect 3516 321574 3568 321580
rect 3422 294400 3478 294409
rect 3422 294335 3478 294344
rect 3528 280129 3556 321574
rect 3620 308825 3648 349114
rect 523684 345092 523736 345098
rect 523684 345034 523736 345040
rect 59358 336016 59414 336025
rect 59358 335951 59414 335960
rect 59372 335374 59400 335951
rect 59360 335368 59412 335374
rect 59360 335310 59412 335316
rect 523696 329905 523724 345034
rect 523788 343233 523816 357410
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580184 345098 580212 346015
rect 580172 345092 580224 345098
rect 580172 345034 580224 345040
rect 523774 343224 523830 343233
rect 523774 343159 523830 343168
rect 523682 329896 523738 329905
rect 523682 329831 523738 329840
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 59358 321736 59414 321745
rect 59358 321671 59414 321680
rect 59372 321638 59400 321671
rect 580184 321638 580212 322623
rect 59360 321632 59412 321638
rect 59360 321574 59412 321580
rect 523500 321632 523552 321638
rect 523500 321574 523552 321580
rect 580172 321632 580224 321638
rect 580172 321574 580224 321580
rect 523512 316577 523540 321574
rect 523498 316568 523554 316577
rect 523498 316503 523554 316512
rect 579802 310856 579858 310865
rect 579802 310791 579858 310800
rect 579816 310554 579844 310791
rect 523684 310548 523736 310554
rect 523684 310490 523736 310496
rect 579804 310548 579856 310554
rect 579804 310490 579856 310496
rect 3606 308816 3662 308825
rect 3606 308751 3662 308760
rect 59358 307456 59414 307465
rect 59358 307391 59414 307400
rect 59372 306406 59400 307391
rect 3700 306400 3752 306406
rect 3700 306342 3752 306348
rect 59360 306400 59412 306406
rect 59360 306342 59412 306348
rect 3608 292596 3660 292602
rect 3608 292538 3660 292544
rect 3514 280120 3570 280129
rect 3514 280055 3570 280064
rect 3424 278792 3476 278798
rect 3424 278734 3476 278740
rect 3436 237017 3464 278734
rect 3620 251297 3648 292538
rect 3712 265713 3740 306342
rect 523696 303249 523724 310490
rect 523682 303240 523738 303249
rect 523682 303175 523738 303184
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 580184 298178 580212 299095
rect 523224 298172 523276 298178
rect 523224 298114 523276 298120
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 59358 293176 59414 293185
rect 59358 293111 59414 293120
rect 59372 292602 59400 293111
rect 59360 292596 59412 292602
rect 59360 292538 59412 292544
rect 523236 289921 523264 298114
rect 523222 289912 523278 289921
rect 523222 289847 523278 289856
rect 59358 278896 59414 278905
rect 59358 278831 59414 278840
rect 59372 278798 59400 278831
rect 59360 278792 59412 278798
rect 59360 278734 59412 278740
rect 524326 276584 524382 276593
rect 524326 276519 524382 276528
rect 524340 276010 524368 276519
rect 524328 276004 524380 276010
rect 524328 275946 524380 275952
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 3698 265704 3754 265713
rect 3698 265639 3754 265648
rect 59358 264616 59414 264625
rect 59358 264551 59414 264560
rect 59372 263634 59400 264551
rect 579802 263936 579858 263945
rect 579802 263871 579858 263880
rect 579816 263634 579844 263871
rect 3700 263628 3752 263634
rect 3700 263570 3752 263576
rect 59360 263628 59412 263634
rect 59360 263570 59412 263576
rect 524328 263628 524380 263634
rect 524328 263570 524380 263576
rect 579804 263628 579856 263634
rect 579804 263570 579856 263576
rect 3606 251288 3662 251297
rect 3606 251223 3662 251232
rect 3516 249824 3568 249830
rect 3516 249766 3568 249772
rect 3422 237008 3478 237017
rect 3422 236943 3478 236952
rect 3424 220856 3476 220862
rect 3424 220798 3476 220804
rect 3436 179489 3464 220798
rect 3528 208185 3556 249766
rect 3608 236020 3660 236026
rect 3608 235962 3660 235968
rect 3514 208176 3570 208185
rect 3514 208111 3570 208120
rect 3620 193905 3648 235962
rect 3712 222601 3740 263570
rect 524340 263265 524368 263570
rect 524326 263256 524382 263265
rect 524326 263191 524382 263200
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 580184 251258 580212 252175
rect 523960 251252 524012 251258
rect 523960 251194 524012 251200
rect 580172 251252 580224 251258
rect 580172 251194 580224 251200
rect 59358 250336 59414 250345
rect 59358 250271 59414 250280
rect 59372 249830 59400 250271
rect 523972 249937 524000 251194
rect 523958 249928 524014 249937
rect 523958 249863 524014 249872
rect 59360 249824 59412 249830
rect 59360 249766 59412 249772
rect 523682 236600 523738 236609
rect 523682 236535 523738 236544
rect 59358 236056 59414 236065
rect 59358 235991 59360 236000
rect 59412 235991 59414 236000
rect 59360 235962 59412 235968
rect 523696 229090 523724 236535
rect 523684 229084 523736 229090
rect 523684 229026 523736 229032
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 523682 223272 523738 223281
rect 523682 223207 523738 223216
rect 3698 222592 3754 222601
rect 3698 222527 3754 222536
rect 59358 221776 59414 221785
rect 59358 221711 59414 221720
rect 59372 220862 59400 221711
rect 59360 220856 59412 220862
rect 59360 220798 59412 220804
rect 523696 218006 523724 223207
rect 523684 218000 523736 218006
rect 523684 217942 523736 217948
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 523406 209944 523462 209953
rect 523406 209879 523462 209888
rect 59358 207496 59414 207505
rect 59358 207431 59414 207440
rect 59372 207058 59400 207431
rect 3700 207052 3752 207058
rect 3700 206994 3752 207000
rect 59360 207052 59412 207058
rect 59360 206994 59412 207000
rect 3606 193896 3662 193905
rect 3606 193831 3662 193840
rect 3608 191888 3660 191894
rect 3608 191830 3660 191836
rect 3422 179480 3478 179489
rect 3422 179415 3478 179424
rect 3516 178084 3568 178090
rect 3516 178026 3568 178032
rect 3424 164280 3476 164286
rect 3424 164222 3476 164228
rect 3436 122097 3464 164222
rect 3528 136377 3556 178026
rect 3620 150793 3648 191830
rect 3712 165073 3740 206994
rect 523420 205630 523448 209879
rect 523408 205624 523460 205630
rect 523408 205566 523460 205572
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 523682 196616 523738 196625
rect 523682 196551 523738 196560
rect 59358 193216 59414 193225
rect 59358 193151 59414 193160
rect 59372 191894 59400 193151
rect 59360 191888 59412 191894
rect 59360 191830 59412 191836
rect 523696 182170 523724 196551
rect 523774 183288 523830 183297
rect 523774 183223 523830 183232
rect 523684 182164 523736 182170
rect 523684 182106 523736 182112
rect 59358 178936 59414 178945
rect 59358 178871 59414 178880
rect 59372 178090 59400 178871
rect 59360 178084 59412 178090
rect 59360 178026 59412 178032
rect 523788 171086 523816 183223
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 523776 171080 523828 171086
rect 523776 171022 523828 171028
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 523682 169960 523738 169969
rect 523682 169895 523738 169904
rect 3698 165064 3754 165073
rect 3698 164999 3754 165008
rect 59358 164656 59414 164665
rect 59358 164591 59414 164600
rect 59372 164286 59400 164591
rect 59360 164280 59412 164286
rect 59360 164222 59412 164228
rect 523696 158710 523724 169895
rect 523684 158704 523736 158710
rect 523684 158646 523736 158652
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 523682 156632 523738 156641
rect 523682 156567 523738 156576
rect 3606 150784 3662 150793
rect 3606 150719 3662 150728
rect 59358 150376 59414 150385
rect 59358 150311 59414 150320
rect 59372 149122 59400 150311
rect 3700 149116 3752 149122
rect 3700 149058 3752 149064
rect 59360 149116 59412 149122
rect 59360 149058 59412 149064
rect 3514 136368 3570 136377
rect 3514 136303 3570 136312
rect 3608 135312 3660 135318
rect 3608 135254 3660 135260
rect 3422 122088 3478 122097
rect 3422 122023 3478 122032
rect 3516 121508 3568 121514
rect 3516 121450 3568 121456
rect 3528 78985 3556 121450
rect 3620 93265 3648 135254
rect 3712 107681 3740 149058
rect 59358 136096 59414 136105
rect 59358 136031 59414 136040
rect 59372 135318 59400 136031
rect 59360 135312 59412 135318
rect 59360 135254 59412 135260
rect 523696 135250 523724 156567
rect 523866 143304 523922 143313
rect 523866 143239 523922 143248
rect 523684 135244 523736 135250
rect 523684 135186 523736 135192
rect 523774 129976 523830 129985
rect 523774 129911 523830 129920
rect 59358 121816 59414 121825
rect 59358 121751 59414 121760
rect 59372 121514 59400 121751
rect 59360 121508 59412 121514
rect 59360 121450 59412 121456
rect 523682 116648 523738 116657
rect 523682 116583 523738 116592
rect 3698 107672 3754 107681
rect 3698 107607 3754 107616
rect 59358 107536 59414 107545
rect 59358 107471 59414 107480
rect 59372 106350 59400 107471
rect 3792 106344 3844 106350
rect 3792 106286 3844 106292
rect 59360 106344 59412 106350
rect 59360 106286 59412 106292
rect 3606 93256 3662 93265
rect 3606 93191 3662 93200
rect 3700 92540 3752 92546
rect 3700 92482 3752 92488
rect 3514 78976 3570 78985
rect 3514 78911 3570 78920
rect 3424 78736 3476 78742
rect 3424 78678 3476 78684
rect 2688 40724 2740 40730
rect 2688 40666 2740 40672
rect 2700 3534 2728 40666
rect 3436 35873 3464 78678
rect 3608 63572 3660 63578
rect 3608 63514 3660 63520
rect 3516 49768 3568 49774
rect 3516 49710 3568 49716
rect 3422 35864 3478 35873
rect 3422 35799 3478 35808
rect 3528 7177 3556 49710
rect 3620 21457 3648 63514
rect 3712 50153 3740 92482
rect 3804 64569 3832 106286
rect 59358 93256 59414 93265
rect 59358 93191 59414 93200
rect 59372 92546 59400 93191
rect 59360 92540 59412 92546
rect 59360 92482 59412 92488
rect 523696 88330 523724 116583
rect 523788 111790 523816 129911
rect 523880 124166 523908 143239
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 523868 124160 523920 124166
rect 523868 124102 523920 124108
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 523776 111784 523828 111790
rect 523776 111726 523828 111732
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 523774 103320 523830 103329
rect 523774 103255 523830 103264
rect 523684 88324 523736 88330
rect 523684 88266 523736 88272
rect 59358 78976 59414 78985
rect 59358 78911 59414 78920
rect 59372 78742 59400 78911
rect 59360 78736 59412 78742
rect 59360 78678 59412 78684
rect 523788 77246 523816 103255
rect 523866 89992 523922 90001
rect 523866 89927 523922 89936
rect 523776 77240 523828 77246
rect 523776 77182 523828 77188
rect 523682 76664 523738 76673
rect 523682 76599 523738 76608
rect 59358 64696 59414 64705
rect 59358 64631 59414 64640
rect 3790 64560 3846 64569
rect 3790 64495 3846 64504
rect 59372 63578 59400 64631
rect 59360 63572 59412 63578
rect 59360 63514 59412 63520
rect 59358 50416 59414 50425
rect 59358 50351 59414 50360
rect 3698 50144 3754 50153
rect 3698 50079 3754 50088
rect 59372 49774 59400 50351
rect 59360 49768 59412 49774
rect 59360 49710 59412 49716
rect 383134 43438 383516 43466
rect 62132 43302 62606 43330
rect 3606 21448 3662 21457
rect 3606 21383 3662 21392
rect 3514 7168 3570 7177
rect 3514 7103 3570 7112
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 62132 3466 62160 43302
rect 63696 40730 63724 43316
rect 63684 40724 63736 40730
rect 63684 40666 63736 40672
rect 64892 40186 64920 43316
rect 64880 40180 64932 40186
rect 64880 40122 64932 40128
rect 66088 40118 66116 43316
rect 67284 40730 67312 43316
rect 68494 43302 68968 43330
rect 69690 43302 70348 43330
rect 67272 40724 67324 40730
rect 67272 40666 67324 40672
rect 66168 40180 66220 40186
rect 66168 40122 66220 40128
rect 66076 40112 66128 40118
rect 66076 40054 66128 40060
rect 66180 4894 66208 40122
rect 66904 40112 66956 40118
rect 66904 40054 66956 40060
rect 66916 15910 66944 40054
rect 66904 15904 66956 15910
rect 66904 15846 66956 15852
rect 66168 4888 66220 4894
rect 66168 4830 66220 4836
rect 68940 4826 68968 43302
rect 70320 17338 70348 43302
rect 70872 40118 70900 43316
rect 72068 40118 72096 43316
rect 70860 40112 70912 40118
rect 70860 40054 70912 40060
rect 71688 40112 71740 40118
rect 71688 40054 71740 40060
rect 72056 40112 72108 40118
rect 72056 40054 72108 40060
rect 73068 40112 73120 40118
rect 73068 40054 73120 40060
rect 70308 17332 70360 17338
rect 70308 17274 70360 17280
rect 68928 4820 68980 4826
rect 68928 4762 68980 4768
rect 71700 3670 71728 40054
rect 73080 18630 73108 40054
rect 73264 39438 73292 43316
rect 74368 43302 74474 43330
rect 75670 43302 75868 43330
rect 73252 39432 73304 39438
rect 73252 39374 73304 39380
rect 73068 18624 73120 18630
rect 73068 18566 73120 18572
rect 71688 3664 71740 3670
rect 71688 3606 71740 3612
rect 74368 3534 74396 43302
rect 75840 19990 75868 43302
rect 76852 37942 76880 43316
rect 78062 43302 78628 43330
rect 79258 43302 80008 43330
rect 76840 37936 76892 37942
rect 76840 37878 76892 37884
rect 75828 19984 75880 19990
rect 75828 19926 75880 19932
rect 78600 3602 78628 43302
rect 79980 21418 80008 43302
rect 80440 40118 80468 43316
rect 81636 41002 81664 43316
rect 81624 40996 81676 41002
rect 81624 40938 81676 40944
rect 82832 40118 82860 43316
rect 84042 43302 84148 43330
rect 85238 43302 85528 43330
rect 86434 43302 86908 43330
rect 87630 43302 88288 43330
rect 80428 40112 80480 40118
rect 80428 40054 80480 40060
rect 81348 40112 81400 40118
rect 81348 40054 81400 40060
rect 82820 40112 82872 40118
rect 82820 40054 82872 40060
rect 84016 40112 84068 40118
rect 84016 40054 84068 40060
rect 79968 21412 80020 21418
rect 79968 21354 80020 21360
rect 81360 14550 81388 40054
rect 84028 22778 84056 40054
rect 84016 22772 84068 22778
rect 84016 22714 84068 22720
rect 81348 14544 81400 14550
rect 81348 14486 81400 14492
rect 84120 13190 84148 43302
rect 84108 13184 84160 13190
rect 84108 13126 84160 13132
rect 78588 3596 78640 3602
rect 78588 3538 78640 3544
rect 74356 3528 74408 3534
rect 85500 3505 85528 43302
rect 86880 24138 86908 43302
rect 86868 24132 86920 24138
rect 86868 24074 86920 24080
rect 88260 3942 88288 43302
rect 88720 40798 88748 43316
rect 88708 40792 88760 40798
rect 88708 40734 88760 40740
rect 89916 40118 89944 43316
rect 91112 40118 91140 43316
rect 89904 40112 89956 40118
rect 89904 40054 89956 40060
rect 91008 40112 91060 40118
rect 91008 40054 91060 40060
rect 91100 40112 91152 40118
rect 91100 40054 91152 40060
rect 91020 25566 91048 40054
rect 91008 25560 91060 25566
rect 91008 25502 91060 25508
rect 88248 3936 88300 3942
rect 88248 3878 88300 3884
rect 74356 3470 74408 3476
rect 85486 3496 85542 3505
rect 62120 3460 62172 3466
rect 85486 3431 85542 3440
rect 62120 3402 62172 3408
rect 92308 3369 92336 43316
rect 93518 43302 93808 43330
rect 94714 43302 95188 43330
rect 92388 40112 92440 40118
rect 92388 40054 92440 40060
rect 92294 3360 92350 3369
rect 92294 3295 92350 3304
rect 92400 3126 92428 40054
rect 93780 26926 93808 43302
rect 93768 26920 93820 26926
rect 93768 26862 93820 26868
rect 95160 3466 95188 43302
rect 95896 40866 95924 43316
rect 95884 40860 95936 40866
rect 95884 40802 95936 40808
rect 97092 40118 97120 43316
rect 98288 40118 98316 43316
rect 99484 40118 99512 43316
rect 100588 43302 100694 43330
rect 101890 43302 102088 43330
rect 97080 40112 97132 40118
rect 97080 40054 97132 40060
rect 97908 40112 97960 40118
rect 97908 40054 97960 40060
rect 98276 40112 98328 40118
rect 98276 40054 98328 40060
rect 99288 40112 99340 40118
rect 99288 40054 99340 40060
rect 99472 40112 99524 40118
rect 99472 40054 99524 40060
rect 97920 28286 97948 40054
rect 97908 28280 97960 28286
rect 97908 28222 97960 28228
rect 95148 3460 95200 3466
rect 95148 3402 95200 3408
rect 92388 3120 92440 3126
rect 92388 3062 92440 3068
rect 99300 3058 99328 40054
rect 100588 6186 100616 43302
rect 100668 40112 100720 40118
rect 100668 40054 100720 40060
rect 100576 6180 100628 6186
rect 100576 6122 100628 6128
rect 100680 3262 100708 40054
rect 102060 29714 102088 43302
rect 103072 40934 103100 43316
rect 104282 43302 104848 43330
rect 103060 40928 103112 40934
rect 103060 40870 103112 40876
rect 102048 29708 102100 29714
rect 102048 29650 102100 29656
rect 104820 7614 104848 43302
rect 105464 40118 105492 43316
rect 106660 40118 106688 43316
rect 107856 40118 107884 43316
rect 109052 40118 109080 43316
rect 110248 41138 110276 43316
rect 111458 43302 111748 43330
rect 112654 43302 113128 43330
rect 110236 41132 110288 41138
rect 110236 41074 110288 41080
rect 105452 40112 105504 40118
rect 105452 40054 105504 40060
rect 106188 40112 106240 40118
rect 106188 40054 106240 40060
rect 106648 40112 106700 40118
rect 106648 40054 106700 40060
rect 107568 40112 107620 40118
rect 107568 40054 107620 40060
rect 107844 40112 107896 40118
rect 107844 40054 107896 40060
rect 108948 40112 109000 40118
rect 108948 40054 109000 40060
rect 109040 40112 109092 40118
rect 109040 40054 109092 40060
rect 110328 40112 110380 40118
rect 110328 40054 110380 40060
rect 106200 31142 106228 40054
rect 106188 31136 106240 31142
rect 106188 31078 106240 31084
rect 104808 7608 104860 7614
rect 104808 7550 104860 7556
rect 100668 3256 100720 3262
rect 100668 3198 100720 3204
rect 107580 3194 107608 40054
rect 108960 8974 108988 40054
rect 110340 32434 110368 40054
rect 110328 32428 110380 32434
rect 110328 32370 110380 32376
rect 111720 10334 111748 43302
rect 113100 33862 113128 43302
rect 113744 40118 113772 43316
rect 114940 40118 114968 43316
rect 116136 40118 116164 43316
rect 117332 40118 117360 43316
rect 113732 40112 113784 40118
rect 113732 40054 113784 40060
rect 114468 40112 114520 40118
rect 114468 40054 114520 40060
rect 114928 40112 114980 40118
rect 114928 40054 114980 40060
rect 115848 40112 115900 40118
rect 115848 40054 115900 40060
rect 116124 40112 116176 40118
rect 116124 40054 116176 40060
rect 117228 40112 117280 40118
rect 117228 40054 117280 40060
rect 117320 40112 117372 40118
rect 117320 40054 117372 40060
rect 113088 33856 113140 33862
rect 113088 33798 113140 33804
rect 111708 10328 111760 10334
rect 111708 10270 111760 10276
rect 108948 8968 109000 8974
rect 108948 8910 109000 8916
rect 114480 3806 114508 40054
rect 115860 11762 115888 40054
rect 117240 35290 117268 40054
rect 117228 35284 117280 35290
rect 117228 35226 117280 35232
rect 118528 13122 118556 43316
rect 118608 40112 118660 40118
rect 118608 40054 118660 40060
rect 118516 13116 118568 13122
rect 118516 13058 118568 13064
rect 115848 11756 115900 11762
rect 115848 11698 115900 11704
rect 118620 4146 118648 40054
rect 119724 36582 119752 43316
rect 120934 43302 121408 43330
rect 122130 43302 122788 43330
rect 119712 36576 119764 36582
rect 119712 36518 119764 36524
rect 118608 4140 118660 4146
rect 118608 4082 118660 4088
rect 114468 3800 114520 3806
rect 114468 3742 114520 3748
rect 121380 3738 121408 43302
rect 122760 14482 122788 43302
rect 123312 38010 123340 43316
rect 124508 40118 124536 43316
rect 125704 40118 125732 43316
rect 124496 40112 124548 40118
rect 124496 40054 124548 40060
rect 125508 40112 125560 40118
rect 125508 40054 125560 40060
rect 125692 40112 125744 40118
rect 125692 40054 125744 40060
rect 126796 40112 126848 40118
rect 126796 40054 126848 40060
rect 123300 38004 123352 38010
rect 123300 37946 123352 37952
rect 122748 14476 122800 14482
rect 122748 14418 122800 14424
rect 121368 3732 121420 3738
rect 121368 3674 121420 3680
rect 125520 3398 125548 40054
rect 126808 15978 126836 40054
rect 126900 39370 126928 43316
rect 128110 43302 128308 43330
rect 129306 43302 129688 43330
rect 130502 43302 131068 43330
rect 126888 39364 126940 39370
rect 126888 39306 126940 39312
rect 126796 15972 126848 15978
rect 126796 15914 126848 15920
rect 126980 15904 127032 15910
rect 126980 15846 127032 15852
rect 126612 4888 126664 4894
rect 126612 4830 126664 4836
rect 125508 3392 125560 3398
rect 125508 3334 125560 3340
rect 107568 3188 107620 3194
rect 107568 3130 107620 3136
rect 99288 3052 99340 3058
rect 99288 2994 99340 3000
rect 126624 480 126652 4830
rect 126992 3482 127020 15846
rect 128280 3874 128308 43302
rect 128452 40724 128504 40730
rect 128452 40666 128504 40672
rect 128268 3868 128320 3874
rect 128268 3810 128320 3816
rect 128464 3482 128492 40666
rect 129660 17270 129688 43302
rect 131040 29782 131068 43302
rect 131684 41070 131712 43316
rect 131672 41064 131724 41070
rect 131672 41006 131724 41012
rect 132880 40118 132908 43316
rect 134076 40118 134104 43316
rect 135272 40118 135300 43316
rect 132868 40112 132920 40118
rect 132868 40054 132920 40060
rect 133788 40112 133840 40118
rect 133788 40054 133840 40060
rect 134064 40112 134116 40118
rect 134064 40054 134116 40060
rect 135168 40112 135220 40118
rect 135168 40054 135220 40060
rect 135260 40112 135312 40118
rect 135260 40054 135312 40060
rect 131028 29776 131080 29782
rect 131028 29718 131080 29724
rect 132592 18624 132644 18630
rect 132592 18566 132644 18572
rect 131120 17332 131172 17338
rect 131120 17274 131172 17280
rect 129648 17264 129700 17270
rect 129648 17206 129700 17212
rect 130200 4820 130252 4826
rect 130200 4762 130252 4768
rect 126992 3454 127848 3482
rect 128464 3454 129044 3482
rect 127820 480 127848 3454
rect 129016 480 129044 3454
rect 130212 480 130240 4762
rect 131132 3482 131160 17274
rect 132500 3664 132552 3670
rect 132500 3606 132552 3612
rect 131132 3454 131436 3482
rect 131408 480 131436 3454
rect 132512 3346 132540 3606
rect 132604 3534 132632 18566
rect 133800 4962 133828 40054
rect 133880 39432 133932 39438
rect 133880 39374 133932 39380
rect 133788 4956 133840 4962
rect 133788 4898 133840 4904
rect 132592 3528 132644 3534
rect 132592 3470 132644 3476
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 132512 3318 132632 3346
rect 132604 480 132632 3318
rect 133800 480 133828 3470
rect 133892 3346 133920 39374
rect 135180 31210 135208 40054
rect 135168 31204 135220 31210
rect 135168 31146 135220 31152
rect 136468 18630 136496 43316
rect 137678 43302 137968 43330
rect 136548 40112 136600 40118
rect 136548 40054 136600 40060
rect 136456 18624 136508 18630
rect 136456 18566 136508 18572
rect 133892 3318 134932 3346
rect 136560 3330 136588 40054
rect 136640 19984 136692 19990
rect 136640 19926 136692 19932
rect 136652 3346 136680 19926
rect 137940 7682 137968 43302
rect 138860 40730 138888 43316
rect 139978 43302 140728 43330
rect 138848 40724 138900 40730
rect 138848 40666 138900 40672
rect 138020 37936 138072 37942
rect 138020 37878 138072 37884
rect 137928 7676 137980 7682
rect 137928 7618 137980 7624
rect 138032 3346 138060 37878
rect 140700 19990 140728 43302
rect 141160 40118 141188 43316
rect 142252 40996 142304 41002
rect 142252 40938 142304 40944
rect 141148 40112 141200 40118
rect 141148 40054 141200 40060
rect 142068 40112 142120 40118
rect 142068 40054 142120 40060
rect 142080 32502 142108 40054
rect 142068 32496 142120 32502
rect 142068 32438 142120 32444
rect 140780 21412 140832 21418
rect 140780 21354 140832 21360
rect 140688 19984 140740 19990
rect 140688 19926 140740 19932
rect 139676 3596 139728 3602
rect 139676 3538 139728 3544
rect 134904 480 134932 3318
rect 136088 3324 136140 3330
rect 136088 3266 136140 3272
rect 136548 3324 136600 3330
rect 136652 3318 137324 3346
rect 138032 3318 138520 3346
rect 136548 3266 136600 3272
rect 136100 480 136128 3266
rect 137296 480 137324 3318
rect 138492 480 138520 3318
rect 139688 480 139716 3538
rect 140792 3482 140820 21354
rect 140872 14544 140924 14550
rect 140872 14486 140924 14492
rect 140884 3602 140912 14486
rect 140872 3596 140924 3602
rect 140872 3538 140924 3544
rect 142068 3596 142120 3602
rect 142068 3538 142120 3544
rect 140792 3454 140912 3482
rect 140884 480 140912 3454
rect 142080 480 142108 3538
rect 142264 3346 142292 40938
rect 142356 40118 142384 43316
rect 143552 40118 143580 43316
rect 142344 40112 142396 40118
rect 142344 40054 142396 40060
rect 143448 40112 143500 40118
rect 143448 40054 143500 40060
rect 143540 40112 143592 40118
rect 143540 40054 143592 40060
rect 143460 4010 143488 40054
rect 144748 33794 144776 43316
rect 145944 41206 145972 43316
rect 147154 43302 147628 43330
rect 148350 43302 149008 43330
rect 145932 41200 145984 41206
rect 145932 41142 145984 41148
rect 144828 40112 144880 40118
rect 144828 40054 144880 40060
rect 144736 33788 144788 33794
rect 144736 33730 144788 33736
rect 143540 22772 143592 22778
rect 143540 22714 143592 22720
rect 143448 4004 143500 4010
rect 143448 3946 143500 3952
rect 143552 3346 143580 22714
rect 144840 21418 144868 40054
rect 147600 22778 147628 43302
rect 148980 35222 149008 43302
rect 149532 40118 149560 43316
rect 150624 40792 150676 40798
rect 150624 40734 150676 40740
rect 149520 40112 149572 40118
rect 149520 40054 149572 40060
rect 150348 40112 150400 40118
rect 150348 40054 150400 40060
rect 148968 35216 149020 35222
rect 148968 35158 149020 35164
rect 147680 24132 147732 24138
rect 147680 24074 147732 24080
rect 147588 22772 147640 22778
rect 147588 22714 147640 22720
rect 144828 21412 144880 21418
rect 144828 21354 144880 21360
rect 144920 13184 144972 13190
rect 144920 13126 144972 13132
rect 144932 3346 144960 13126
rect 146850 3496 146906 3505
rect 146850 3431 146906 3440
rect 142264 3318 143304 3346
rect 143552 3318 144500 3346
rect 144932 3318 145696 3346
rect 143276 480 143304 3318
rect 144472 480 144500 3318
rect 145668 480 145696 3318
rect 146864 480 146892 3431
rect 147692 3346 147720 24074
rect 150360 4078 150388 40054
rect 150532 25560 150584 25566
rect 150532 25502 150584 25508
rect 150348 4072 150400 4078
rect 150348 4014 150400 4020
rect 149244 3936 149296 3942
rect 149244 3878 149296 3884
rect 147692 3318 148088 3346
rect 148060 480 148088 3318
rect 149256 480 149284 3878
rect 150544 3602 150572 25502
rect 150532 3596 150584 3602
rect 150532 3538 150584 3544
rect 150636 3482 150664 40734
rect 150728 40118 150756 43316
rect 150716 40112 150768 40118
rect 150716 40054 150768 40060
rect 151728 40112 151780 40118
rect 151728 40054 151780 40060
rect 151740 24138 151768 40054
rect 151924 36650 151952 43316
rect 151912 36644 151964 36650
rect 151912 36586 151964 36592
rect 151728 24132 151780 24138
rect 151728 24074 151780 24080
rect 153120 3670 153148 43316
rect 154330 43302 154528 43330
rect 154500 25566 154528 43302
rect 155512 37942 155540 43316
rect 156722 43302 157288 43330
rect 155500 37936 155552 37942
rect 155500 37878 155552 37884
rect 154580 26920 154632 26926
rect 154580 26862 154632 26868
rect 154488 25560 154540 25566
rect 154488 25502 154540 25508
rect 153108 3664 153160 3670
rect 153108 3606 153160 3612
rect 151544 3596 151596 3602
rect 151544 3538 151596 3544
rect 150452 3454 150664 3482
rect 150452 480 150480 3454
rect 151556 480 151584 3538
rect 153934 3360 153990 3369
rect 154592 3346 154620 26862
rect 157260 3602 157288 43302
rect 157432 40860 157484 40866
rect 157432 40802 157484 40808
rect 157248 3596 157300 3602
rect 157248 3538 157300 3544
rect 156328 3460 156380 3466
rect 156328 3402 156380 3408
rect 154592 3318 155172 3346
rect 153934 3295 153990 3304
rect 152740 3120 152792 3126
rect 152740 3062 152792 3068
rect 152752 480 152780 3062
rect 153948 480 153976 3295
rect 155144 480 155172 3318
rect 156340 480 156368 3402
rect 157444 1578 157472 40802
rect 157904 40118 157932 43316
rect 157892 40112 157944 40118
rect 157892 40054 157944 40060
rect 158628 40112 158680 40118
rect 158628 40054 158680 40060
rect 158640 26926 158668 40054
rect 159100 39438 159128 43316
rect 160296 40118 160324 43316
rect 161492 40118 161520 43316
rect 160284 40112 160336 40118
rect 160284 40054 160336 40060
rect 161388 40112 161440 40118
rect 161388 40054 161440 40060
rect 161480 40112 161532 40118
rect 161480 40054 161532 40060
rect 159088 39432 159140 39438
rect 159088 39374 159140 39380
rect 158812 28280 158864 28286
rect 158812 28222 158864 28228
rect 158628 26920 158680 26926
rect 158628 26862 158680 26868
rect 158824 1578 158852 28222
rect 161400 3942 161428 40054
rect 162688 29646 162716 43316
rect 163898 43302 164188 43330
rect 165002 43302 165568 43330
rect 162768 40112 162820 40118
rect 162768 40054 162820 40060
rect 162676 29640 162728 29646
rect 162676 29582 162728 29588
rect 162780 6322 162808 40054
rect 162860 29708 162912 29714
rect 162860 29650 162912 29656
rect 162768 6316 162820 6322
rect 162768 6258 162820 6264
rect 162308 6180 162360 6186
rect 162308 6122 162360 6128
rect 161388 3936 161440 3942
rect 161388 3878 161440 3884
rect 161112 3256 161164 3262
rect 161112 3198 161164 3204
rect 159916 3052 159968 3058
rect 159916 2994 159968 3000
rect 157444 1550 157564 1578
rect 157536 480 157564 1550
rect 158732 1550 158852 1578
rect 158732 480 158760 1550
rect 159928 480 159956 2994
rect 161124 480 161152 3198
rect 162320 480 162348 6122
rect 162872 3482 162900 29650
rect 162872 3454 163544 3482
rect 164160 3466 164188 43302
rect 164332 40928 164384 40934
rect 164332 40870 164384 40876
rect 164344 3482 164372 40870
rect 165540 28286 165568 43302
rect 166184 40118 166212 43316
rect 167380 41206 167408 43316
rect 167368 41200 167420 41206
rect 167368 41142 167420 41148
rect 168576 40118 168604 43316
rect 169772 40118 169800 43316
rect 170982 43302 171088 43330
rect 172178 43302 172468 43330
rect 173374 43302 173848 43330
rect 166172 40112 166224 40118
rect 166172 40054 166224 40060
rect 166908 40112 166960 40118
rect 166908 40054 166960 40060
rect 168564 40112 168616 40118
rect 168564 40054 168616 40060
rect 169668 40112 169720 40118
rect 169668 40054 169720 40060
rect 169760 40112 169812 40118
rect 169760 40054 169812 40060
rect 170956 40112 171008 40118
rect 170956 40054 171008 40060
rect 166920 31074 166948 40054
rect 167092 31136 167144 31142
rect 167092 31078 167144 31084
rect 166908 31068 166960 31074
rect 166908 31010 166960 31016
rect 165528 28280 165580 28286
rect 165528 28222 165580 28228
rect 165896 7608 165948 7614
rect 165896 7550 165948 7556
rect 163516 480 163544 3454
rect 164148 3460 164200 3466
rect 164344 3454 164740 3482
rect 164148 3402 164200 3408
rect 164712 480 164740 3454
rect 165908 480 165936 7550
rect 167104 480 167132 31078
rect 169392 8968 169444 8974
rect 169392 8910 169444 8916
rect 168196 3188 168248 3194
rect 168196 3130 168248 3136
rect 168208 480 168236 3130
rect 169404 480 169432 8910
rect 169680 7614 169708 40054
rect 170968 32434 170996 40054
rect 169760 32428 169812 32434
rect 169760 32370 169812 32376
rect 170956 32428 171008 32434
rect 170956 32370 171008 32376
rect 169668 7608 169720 7614
rect 169668 7550 169720 7556
rect 169772 3482 169800 32370
rect 171060 3534 171088 43302
rect 171232 41132 171284 41138
rect 171232 41074 171284 41080
rect 171048 3528 171100 3534
rect 169772 3454 170628 3482
rect 171048 3470 171100 3476
rect 170600 480 170628 3454
rect 171244 3346 171272 41074
rect 172440 8974 172468 43302
rect 172520 10328 172572 10334
rect 172520 10270 172572 10276
rect 172428 8968 172480 8974
rect 172428 8910 172480 8916
rect 172532 3346 172560 10270
rect 173820 4826 173848 43302
rect 174556 40934 174584 43316
rect 174544 40928 174596 40934
rect 174544 40870 174596 40876
rect 175752 40118 175780 43316
rect 176948 40118 176976 43316
rect 178144 40118 178172 43316
rect 179248 43302 179354 43330
rect 180550 43302 180748 43330
rect 175740 40112 175792 40118
rect 175740 40054 175792 40060
rect 176568 40112 176620 40118
rect 176568 40054 176620 40060
rect 176936 40112 176988 40118
rect 176936 40054 176988 40060
rect 177948 40112 178000 40118
rect 177948 40054 178000 40060
rect 178132 40112 178184 40118
rect 178132 40054 178184 40060
rect 173900 33856 173952 33862
rect 173900 33798 173952 33804
rect 173808 4820 173860 4826
rect 173808 4762 173860 4768
rect 173912 3346 173940 33798
rect 175372 11756 175424 11762
rect 175372 11698 175424 11704
rect 175280 3800 175332 3806
rect 175280 3742 175332 3748
rect 171244 3318 171824 3346
rect 172532 3318 173020 3346
rect 173912 3318 174216 3346
rect 171796 480 171824 3318
rect 172992 480 173020 3318
rect 174188 480 174216 3318
rect 175292 3074 175320 3742
rect 175384 3262 175412 11698
rect 176580 10402 176608 40054
rect 176660 35284 176712 35290
rect 176660 35226 176712 35232
rect 176568 10396 176620 10402
rect 176568 10338 176620 10344
rect 176672 3346 176700 35226
rect 177960 33930 177988 40054
rect 177948 33924 178000 33930
rect 177948 33866 178000 33872
rect 179248 11762 179276 43302
rect 179328 40112 179380 40118
rect 179328 40054 179380 40060
rect 179236 11756 179288 11762
rect 179236 11698 179288 11704
rect 179340 4146 179368 40054
rect 180720 35290 180748 43302
rect 181732 40866 181760 43316
rect 182942 43302 183508 43330
rect 181720 40860 181772 40866
rect 181720 40802 181772 40808
rect 180800 36576 180852 36582
rect 180800 36518 180852 36524
rect 180708 35284 180760 35290
rect 180708 35226 180760 35232
rect 179420 13116 179472 13122
rect 179420 13058 179472 13064
rect 178960 4140 179012 4146
rect 178960 4082 179012 4088
rect 179328 4140 179380 4146
rect 179328 4082 179380 4088
rect 176672 3318 177804 3346
rect 175372 3256 175424 3262
rect 175372 3198 175424 3204
rect 176568 3256 176620 3262
rect 176568 3198 176620 3204
rect 175292 3046 175412 3074
rect 175384 480 175412 3046
rect 176580 480 176608 3198
rect 177776 480 177804 3318
rect 178972 480 179000 4082
rect 179432 3346 179460 13058
rect 180812 3346 180840 36518
rect 183480 13122 183508 43302
rect 183560 38004 183612 38010
rect 183560 37946 183612 37952
rect 183468 13116 183520 13122
rect 183468 13058 183520 13064
rect 182548 3732 182600 3738
rect 182548 3674 182600 3680
rect 179432 3318 180196 3346
rect 180812 3318 181392 3346
rect 180168 480 180196 3318
rect 181364 480 181392 3318
rect 182560 480 182588 3674
rect 183572 3398 183600 37946
rect 184124 36718 184152 43316
rect 185320 40118 185348 43316
rect 186516 40118 186544 43316
rect 187726 43302 188016 43330
rect 185308 40112 185360 40118
rect 185308 40054 185360 40060
rect 186228 40112 186280 40118
rect 186228 40054 186280 40060
rect 186504 40112 186556 40118
rect 186504 40054 186556 40060
rect 187608 40112 187660 40118
rect 187608 40054 187660 40060
rect 184112 36712 184164 36718
rect 184112 36654 184164 36660
rect 183652 14476 183704 14482
rect 183652 14418 183704 14424
rect 183664 3482 183692 14418
rect 183664 3454 183784 3482
rect 183560 3392 183612 3398
rect 183560 3334 183612 3340
rect 183756 480 183784 3454
rect 184848 3392 184900 3398
rect 184848 3334 184900 3340
rect 184860 480 184888 3334
rect 186044 3256 186096 3262
rect 186044 3198 186096 3204
rect 186056 480 186084 3198
rect 186240 3194 186268 40054
rect 186320 15972 186372 15978
rect 186320 15914 186372 15920
rect 186332 3346 186360 15914
rect 187620 14482 187648 40054
rect 187700 39364 187752 39370
rect 187700 39306 187752 39312
rect 187608 14476 187660 14482
rect 187608 14418 187660 14424
rect 187712 3346 187740 39306
rect 187988 38078 188016 43302
rect 188908 41138 188936 43316
rect 190118 43302 190408 43330
rect 191222 43302 191788 43330
rect 192418 43302 193168 43330
rect 188896 41132 188948 41138
rect 188896 41074 188948 41080
rect 187976 38072 188028 38078
rect 187976 38014 188028 38020
rect 190380 4894 190408 43302
rect 191760 29850 191788 43302
rect 191748 29844 191800 29850
rect 191748 29786 191800 29792
rect 191840 29776 191892 29782
rect 191840 29718 191892 29724
rect 190460 17264 190512 17270
rect 190460 17206 190512 17212
rect 190368 4888 190420 4894
rect 190368 4830 190420 4836
rect 189632 3868 189684 3874
rect 189632 3810 189684 3816
rect 186332 3318 187280 3346
rect 187712 3318 188476 3346
rect 186228 3188 186280 3194
rect 186228 3130 186280 3136
rect 187252 480 187280 3318
rect 188448 480 188476 3318
rect 189644 480 189672 3810
rect 190472 3346 190500 17206
rect 191852 3346 191880 29718
rect 190472 3318 190868 3346
rect 191852 3318 192064 3346
rect 190840 480 190868 3318
rect 192036 480 192064 3318
rect 193140 3262 193168 43302
rect 193404 41064 193456 41070
rect 193404 41006 193456 41012
rect 193416 3346 193444 41006
rect 193600 40118 193628 43316
rect 193588 40112 193640 40118
rect 193588 40054 193640 40060
rect 194508 40112 194560 40118
rect 194508 40054 194560 40060
rect 194520 15910 194548 40054
rect 194796 39370 194824 43316
rect 195992 40118 196020 43316
rect 195980 40112 196032 40118
rect 195980 40054 196032 40060
rect 194784 39364 194836 39370
rect 194784 39306 194836 39312
rect 194600 31204 194652 31210
rect 194600 31146 194652 31152
rect 194508 15904 194560 15910
rect 194508 15846 194560 15852
rect 194416 4956 194468 4962
rect 194416 4898 194468 4904
rect 193232 3318 193444 3346
rect 193128 3256 193180 3262
rect 193128 3198 193180 3204
rect 193232 480 193260 3318
rect 194428 480 194456 4898
rect 194612 3346 194640 31146
rect 197188 17270 197216 43316
rect 198398 43302 198688 43330
rect 199594 43302 200068 43330
rect 200790 43302 201448 43330
rect 197268 40112 197320 40118
rect 197268 40054 197320 40060
rect 197176 17264 197228 17270
rect 197176 17206 197228 17212
rect 197280 3874 197308 40054
rect 198660 31142 198688 43302
rect 198648 31136 198700 31142
rect 198648 31078 198700 31084
rect 197360 18624 197412 18630
rect 197360 18566 197412 18572
rect 197268 3868 197320 3874
rect 197268 3810 197320 3816
rect 197372 3346 197400 18566
rect 199200 7676 199252 7682
rect 199200 7618 199252 7624
rect 194612 3318 195652 3346
rect 195624 480 195652 3318
rect 196808 3324 196860 3330
rect 197372 3318 198044 3346
rect 196808 3266 196860 3272
rect 196820 480 196848 3266
rect 198016 480 198044 3318
rect 199212 480 199240 7618
rect 200040 3806 200068 43302
rect 200212 40724 200264 40730
rect 200212 40666 200264 40672
rect 200028 3800 200080 3806
rect 200028 3742 200080 3748
rect 200224 3346 200252 40666
rect 201420 18630 201448 43302
rect 201972 40118 202000 43316
rect 203168 40118 203196 43316
rect 204364 40118 204392 43316
rect 205468 43302 205574 43330
rect 206770 43302 206968 43330
rect 207966 43302 208348 43330
rect 209162 43302 209728 43330
rect 201960 40112 202012 40118
rect 201960 40054 202012 40060
rect 202788 40112 202840 40118
rect 202788 40054 202840 40060
rect 203156 40112 203208 40118
rect 203156 40054 203208 40060
rect 204168 40112 204220 40118
rect 204168 40054 204220 40060
rect 204352 40112 204404 40118
rect 204352 40054 204404 40060
rect 202800 32502 202828 40054
rect 201500 32496 201552 32502
rect 201500 32438 201552 32444
rect 202788 32496 202840 32502
rect 202788 32438 202840 32444
rect 201408 18624 201460 18630
rect 201408 18566 201460 18572
rect 201512 3738 201540 32438
rect 201592 19984 201644 19990
rect 201592 19926 201644 19932
rect 201500 3732 201552 3738
rect 201500 3674 201552 3680
rect 201604 3482 201632 19926
rect 203892 4004 203944 4010
rect 203892 3946 203944 3952
rect 202696 3732 202748 3738
rect 202696 3674 202748 3680
rect 201512 3454 201632 3482
rect 200224 3318 200436 3346
rect 200408 480 200436 3318
rect 201512 480 201540 3454
rect 202708 480 202736 3674
rect 203904 480 203932 3946
rect 204180 3398 204208 40054
rect 205468 33862 205496 43302
rect 205548 40112 205600 40118
rect 205548 40054 205600 40060
rect 205456 33856 205508 33862
rect 205456 33798 205508 33804
rect 205560 21418 205588 40054
rect 205640 33788 205692 33794
rect 205640 33730 205692 33736
rect 204260 21412 204312 21418
rect 204260 21354 204312 21360
rect 205548 21412 205600 21418
rect 205548 21354 205600 21360
rect 204168 3392 204220 3398
rect 204168 3334 204220 3340
rect 204272 3346 204300 21354
rect 205652 3346 205680 33730
rect 206940 3738 206968 43302
rect 207112 40996 207164 41002
rect 207112 40938 207164 40944
rect 206928 3732 206980 3738
rect 206928 3674 206980 3680
rect 207124 3346 207152 40938
rect 208320 19990 208348 43302
rect 208400 22772 208452 22778
rect 208400 22714 208452 22720
rect 208308 19984 208360 19990
rect 208308 19926 208360 19932
rect 208412 3346 208440 22714
rect 209700 6186 209728 43302
rect 210344 41002 210372 43316
rect 210332 40996 210384 41002
rect 210332 40938 210384 40944
rect 211540 40118 211568 43316
rect 212736 40118 212764 43316
rect 213932 40118 213960 43316
rect 211528 40112 211580 40118
rect 211528 40054 211580 40060
rect 212448 40112 212500 40118
rect 212448 40054 212500 40060
rect 212724 40112 212776 40118
rect 212724 40054 212776 40060
rect 213828 40112 213880 40118
rect 213828 40054 213880 40060
rect 213920 40112 213972 40118
rect 213920 40054 213972 40060
rect 209872 35216 209924 35222
rect 209872 35158 209924 35164
rect 209688 6180 209740 6186
rect 209688 6122 209740 6128
rect 204272 3318 205128 3346
rect 205652 3318 206324 3346
rect 207124 3318 207520 3346
rect 208412 3318 208716 3346
rect 205100 480 205128 3318
rect 206296 480 206324 3318
rect 207492 480 207520 3318
rect 208688 480 208716 3318
rect 209884 480 209912 35158
rect 212460 24138 212488 40054
rect 212540 36644 212592 36650
rect 212540 36586 212592 36592
rect 211160 24132 211212 24138
rect 211160 24074 211212 24080
rect 212448 24132 212500 24138
rect 212448 24074 212500 24080
rect 211068 4072 211120 4078
rect 211068 4014 211120 4020
rect 211080 480 211108 4014
rect 211172 3346 211200 24074
rect 212552 3346 212580 36586
rect 213840 35358 213868 40054
rect 213828 35352 213880 35358
rect 213828 35294 213880 35300
rect 215128 22778 215156 43316
rect 215208 40112 215260 40118
rect 215208 40054 215260 40060
rect 215116 22772 215168 22778
rect 215116 22714 215168 22720
rect 214656 3664 214708 3670
rect 214656 3606 214708 3612
rect 211172 3318 212304 3346
rect 212552 3318 213500 3346
rect 212276 480 212304 3318
rect 213472 480 213500 3318
rect 214668 480 214696 3606
rect 215220 3330 215248 40054
rect 216232 36582 216260 43316
rect 217428 40730 217456 43316
rect 217416 40724 217468 40730
rect 217416 40666 217468 40672
rect 218624 40118 218652 43316
rect 218612 40112 218664 40118
rect 218612 40054 218664 40060
rect 219348 40112 219400 40118
rect 219348 40054 219400 40060
rect 216680 37936 216732 37942
rect 216680 37878 216732 37884
rect 216220 36576 216272 36582
rect 216220 36518 216272 36524
rect 215300 25560 215352 25566
rect 215300 25502 215352 25508
rect 215312 3346 215340 25502
rect 216692 3346 216720 37878
rect 218152 26920 218204 26926
rect 218152 26862 218204 26868
rect 218164 3602 218192 26862
rect 219360 6254 219388 40054
rect 219440 39432 219492 39438
rect 219440 39374 219492 39380
rect 219348 6248 219400 6254
rect 219348 6190 219400 6196
rect 218060 3596 218112 3602
rect 218060 3538 218112 3544
rect 218152 3596 218204 3602
rect 218152 3538 218204 3544
rect 219348 3596 219400 3602
rect 219348 3538 219400 3544
rect 218072 3482 218100 3538
rect 218072 3454 218192 3482
rect 215208 3324 215260 3330
rect 215312 3318 215892 3346
rect 216692 3318 217088 3346
rect 215208 3266 215260 3272
rect 215864 480 215892 3318
rect 217060 480 217088 3318
rect 218164 480 218192 3454
rect 219360 480 219388 3538
rect 219452 3346 219480 39374
rect 219820 38010 219848 43316
rect 221016 40118 221044 43316
rect 222212 40118 222240 43316
rect 221004 40112 221056 40118
rect 221004 40054 221056 40060
rect 222108 40112 222160 40118
rect 222108 40054 222160 40060
rect 222200 40112 222252 40118
rect 222200 40054 222252 40060
rect 219808 38004 219860 38010
rect 219808 37946 219860 37952
rect 221740 3936 221792 3942
rect 221740 3878 221792 3884
rect 219452 3318 220584 3346
rect 220556 480 220584 3318
rect 221752 480 221780 3878
rect 222120 3126 222148 40054
rect 223408 29714 223436 43316
rect 224604 40798 224632 43316
rect 225814 43302 226288 43330
rect 224592 40792 224644 40798
rect 224592 40734 224644 40740
rect 223488 40112 223540 40118
rect 223488 40054 223540 40060
rect 223396 29708 223448 29714
rect 223396 29650 223448 29656
rect 223500 7682 223528 40054
rect 223580 29640 223632 29646
rect 223580 29582 223632 29588
rect 223488 7676 223540 7682
rect 223488 7618 223540 7624
rect 222936 6316 222988 6322
rect 222936 6258 222988 6264
rect 222108 3120 222160 3126
rect 222108 3062 222160 3068
rect 222948 480 222976 6258
rect 223592 3346 223620 29582
rect 226260 25566 226288 43302
rect 226996 39438 227024 43316
rect 227904 41200 227956 41206
rect 227904 41142 227956 41148
rect 226984 39432 227036 39438
rect 226984 39374 227036 39380
rect 227812 31068 227864 31074
rect 227812 31010 227864 31016
rect 226340 28280 226392 28286
rect 226340 28222 226392 28228
rect 226248 25560 226300 25566
rect 226248 25502 226300 25508
rect 225328 3460 225380 3466
rect 225328 3402 225380 3408
rect 223592 3318 224172 3346
rect 224144 480 224172 3318
rect 225340 480 225368 3402
rect 226352 3346 226380 28222
rect 227824 3482 227852 31010
rect 227732 3454 227852 3482
rect 226352 3318 226564 3346
rect 226536 480 226564 3318
rect 227732 480 227760 3454
rect 227916 3346 227944 41142
rect 228192 40118 228220 43316
rect 229388 40118 229416 43316
rect 230584 40118 230612 43316
rect 228180 40112 228232 40118
rect 228180 40054 228232 40060
rect 229008 40112 229060 40118
rect 229008 40054 229060 40060
rect 229376 40112 229428 40118
rect 229376 40054 229428 40060
rect 230388 40112 230440 40118
rect 230388 40054 230440 40060
rect 230572 40112 230624 40118
rect 230572 40054 230624 40060
rect 231676 40112 231728 40118
rect 231676 40054 231728 40060
rect 229020 3942 229048 40054
rect 230400 9042 230428 40054
rect 230480 32428 230532 32434
rect 230480 32370 230532 32376
rect 230388 9036 230440 9042
rect 230388 8978 230440 8984
rect 230112 7608 230164 7614
rect 230112 7550 230164 7556
rect 229008 3936 229060 3942
rect 229008 3878 229060 3884
rect 227916 3318 228956 3346
rect 228928 480 228956 3318
rect 230124 480 230152 7550
rect 230492 3482 230520 32370
rect 231688 31074 231716 40054
rect 231676 31068 231728 31074
rect 231676 31010 231728 31016
rect 231780 4010 231808 43316
rect 232990 43302 233188 43330
rect 234186 43302 234568 43330
rect 235382 43302 235948 43330
rect 236578 43302 237328 43330
rect 233160 10334 233188 43302
rect 234540 32434 234568 43302
rect 234528 32428 234580 32434
rect 234528 32370 234580 32376
rect 233148 10328 233200 10334
rect 233148 10270 233200 10276
rect 233700 8968 233752 8974
rect 233700 8910 233752 8916
rect 231768 4004 231820 4010
rect 231768 3946 231820 3952
rect 232504 3528 232556 3534
rect 230492 3454 231348 3482
rect 232504 3470 232556 3476
rect 231320 480 231348 3454
rect 232516 480 232544 3470
rect 233712 480 233740 8910
rect 234804 4820 234856 4826
rect 234804 4762 234856 4768
rect 234816 480 234844 4762
rect 235920 3670 235948 43302
rect 236184 40928 236236 40934
rect 236184 40870 236236 40876
rect 236092 10396 236144 10402
rect 236092 10338 236144 10344
rect 235908 3664 235960 3670
rect 235908 3606 235960 3612
rect 236104 3602 236132 10338
rect 236092 3596 236144 3602
rect 236092 3538 236144 3544
rect 236196 3482 236224 40870
rect 237300 26926 237328 43302
rect 237760 40118 237788 43316
rect 238956 40118 238984 43316
rect 240152 40118 240180 43316
rect 237748 40112 237800 40118
rect 237748 40054 237800 40060
rect 238668 40112 238720 40118
rect 238668 40054 238720 40060
rect 238944 40112 238996 40118
rect 238944 40054 238996 40060
rect 240048 40112 240100 40118
rect 240048 40054 240100 40060
rect 240140 40112 240192 40118
rect 240140 40054 240192 40060
rect 238680 33930 238708 40054
rect 237380 33924 237432 33930
rect 237380 33866 237432 33872
rect 238668 33924 238720 33930
rect 238668 33866 238720 33872
rect 237288 26920 237340 26926
rect 237288 26862 237340 26868
rect 237196 3596 237248 3602
rect 237196 3538 237248 3544
rect 236012 3454 236224 3482
rect 236012 480 236040 3454
rect 237208 480 237236 3538
rect 237392 3482 237420 33866
rect 239588 4140 239640 4146
rect 239588 4082 239640 4088
rect 237392 3454 238432 3482
rect 238404 480 238432 3454
rect 239600 480 239628 4082
rect 240060 4078 240088 40054
rect 241348 35222 241376 43316
rect 242466 43302 242848 43330
rect 243662 43302 244228 43330
rect 241428 40112 241480 40118
rect 241428 40054 241480 40060
rect 241336 35216 241388 35222
rect 241336 35158 241388 35164
rect 241440 11762 241468 40054
rect 241520 35284 241572 35290
rect 241520 35226 241572 35232
rect 240140 11756 240192 11762
rect 240140 11698 240192 11704
rect 241428 11756 241480 11762
rect 241428 11698 241480 11704
rect 240048 4072 240100 4078
rect 240048 4014 240100 4020
rect 240152 3346 240180 11698
rect 241532 3346 241560 35226
rect 242820 3466 242848 43302
rect 242992 40860 243044 40866
rect 242992 40802 243044 40808
rect 242808 3460 242860 3466
rect 242808 3402 242860 3408
rect 243004 3346 243032 40802
rect 244200 28286 244228 43302
rect 244844 36718 244872 43316
rect 246040 40118 246068 43316
rect 247236 40594 247264 43316
rect 248446 43302 248736 43330
rect 249642 43302 249748 43330
rect 250838 43302 251128 43330
rect 252034 43302 252508 43330
rect 247224 40588 247276 40594
rect 247224 40530 247276 40536
rect 248328 40588 248380 40594
rect 248328 40530 248380 40536
rect 246028 40112 246080 40118
rect 246028 40054 246080 40060
rect 246948 40112 247000 40118
rect 246948 40054 247000 40060
rect 244280 36712 244332 36718
rect 244280 36654 244332 36660
rect 244832 36712 244884 36718
rect 244832 36654 244884 36660
rect 244188 28280 244240 28286
rect 244188 28222 244240 28228
rect 244292 3534 244320 36654
rect 244372 13116 244424 13122
rect 244372 13058 244424 13064
rect 244280 3528 244332 3534
rect 244280 3470 244332 3476
rect 240152 3318 240824 3346
rect 241532 3318 242020 3346
rect 243004 3318 243216 3346
rect 240796 480 240824 3318
rect 241992 480 242020 3318
rect 243188 480 243216 3318
rect 244384 480 244412 13058
rect 246960 4010 246988 40054
rect 247040 14476 247092 14482
rect 247040 14418 247092 14424
rect 246948 4004 247000 4010
rect 246948 3946 247000 3952
rect 245568 3528 245620 3534
rect 245568 3470 245620 3476
rect 245580 480 245608 3470
rect 247052 3346 247080 14418
rect 248340 13190 248368 40530
rect 248420 38072 248472 38078
rect 248420 38014 248472 38020
rect 248328 13184 248380 13190
rect 248328 13126 248380 13132
rect 248432 3346 248460 38014
rect 248708 37942 248736 43302
rect 248696 37936 248748 37942
rect 248696 37878 248748 37884
rect 249720 3534 249748 43302
rect 249892 41132 249944 41138
rect 249892 41074 249944 41080
rect 249708 3528 249760 3534
rect 249708 3470 249760 3476
rect 249904 3346 249932 41074
rect 251100 14482 251128 43302
rect 251088 14476 251140 14482
rect 251088 14418 251140 14424
rect 251456 4888 251508 4894
rect 251456 4830 251508 4836
rect 247052 3318 248000 3346
rect 248432 3318 249196 3346
rect 249904 3318 250392 3346
rect 246764 3188 246816 3194
rect 246764 3130 246816 3136
rect 246776 480 246804 3130
rect 247972 480 248000 3318
rect 249168 480 249196 3318
rect 250364 480 250392 3318
rect 251468 480 251496 4830
rect 252480 4826 252508 43302
rect 253216 41206 253244 43316
rect 253204 41200 253256 41206
rect 253204 41142 253256 41148
rect 254412 40118 254440 43316
rect 255608 40118 255636 43316
rect 256804 40118 256832 43316
rect 257908 43302 258014 43330
rect 254400 40112 254452 40118
rect 254400 40054 254452 40060
rect 255228 40112 255280 40118
rect 255228 40054 255280 40060
rect 255596 40112 255648 40118
rect 255596 40054 255648 40060
rect 256608 40112 256660 40118
rect 256608 40054 256660 40060
rect 256792 40112 256844 40118
rect 256792 40054 256844 40060
rect 252652 29844 252704 29850
rect 252652 29786 252704 29792
rect 252468 4820 252520 4826
rect 252468 4762 252520 4768
rect 252664 480 252692 29786
rect 253940 15904 253992 15910
rect 253940 15846 253992 15852
rect 253952 3346 253980 15846
rect 255240 4962 255268 40054
rect 255320 39364 255372 39370
rect 255320 39306 255372 39312
rect 255228 4956 255280 4962
rect 255228 4898 255280 4904
rect 255332 3346 255360 39306
rect 256620 29782 256648 40054
rect 256608 29776 256660 29782
rect 256608 29718 256660 29724
rect 257908 15910 257936 43302
rect 257988 40112 258040 40118
rect 257988 40054 258040 40060
rect 257896 15904 257948 15910
rect 257896 15846 257948 15852
rect 258000 3874 258028 40054
rect 259196 39370 259224 43316
rect 260392 40866 260420 43316
rect 261602 43302 262168 43330
rect 260380 40860 260432 40866
rect 260380 40802 260432 40808
rect 259184 39364 259236 39370
rect 259184 39306 259236 39312
rect 259460 31136 259512 31142
rect 259460 31078 259512 31084
rect 258080 17264 258132 17270
rect 258080 17206 258132 17212
rect 257436 3868 257488 3874
rect 257436 3810 257488 3816
rect 257988 3868 258040 3874
rect 257988 3810 258040 3816
rect 253952 3318 255084 3346
rect 255332 3318 256280 3346
rect 253848 3256 253900 3262
rect 253848 3198 253900 3204
rect 253860 480 253888 3198
rect 255056 480 255084 3318
rect 256252 480 256280 3318
rect 257448 480 257476 3810
rect 258092 3482 258120 17206
rect 259472 3482 259500 31078
rect 262140 17270 262168 43302
rect 262784 40118 262812 43316
rect 263980 40118 264008 43316
rect 265176 40118 265204 43316
rect 262772 40112 262824 40118
rect 262772 40054 262824 40060
rect 263508 40112 263560 40118
rect 263508 40054 263560 40060
rect 263968 40112 264020 40118
rect 263968 40054 264020 40060
rect 264888 40112 264940 40118
rect 264888 40054 264940 40060
rect 265164 40112 265216 40118
rect 265164 40054 265216 40060
rect 266268 40112 266320 40118
rect 266268 40054 266320 40060
rect 262220 32496 262272 32502
rect 262220 32438 262272 32444
rect 262128 17264 262180 17270
rect 262128 17206 262180 17212
rect 262232 3806 262260 32438
rect 263520 31142 263548 40054
rect 263508 31136 263560 31142
rect 263508 31078 263560 31084
rect 262312 18624 262364 18630
rect 262312 18566 262364 18572
rect 261024 3800 261076 3806
rect 261024 3742 261076 3748
rect 262220 3800 262272 3806
rect 262220 3742 262272 3748
rect 258092 3454 258672 3482
rect 259472 3454 259868 3482
rect 258644 480 258672 3454
rect 259840 480 259868 3454
rect 261036 480 261064 3742
rect 262324 3482 262352 18566
rect 264900 4146 264928 40054
rect 264980 21412 265032 21418
rect 264980 21354 265032 21360
rect 264888 4140 264940 4146
rect 264888 4082 264940 4088
rect 263416 3800 263468 3806
rect 263416 3742 263468 3748
rect 262232 3454 262352 3482
rect 262232 480 262260 3454
rect 263428 480 263456 3742
rect 264992 3482 265020 21354
rect 266280 18630 266308 40054
rect 266372 36938 266400 43316
rect 267490 43302 267688 43330
rect 268686 43302 269068 43330
rect 269882 43302 270448 43330
rect 267660 40934 267688 43302
rect 267648 40928 267700 40934
rect 267648 40870 267700 40876
rect 266372 36910 266584 36938
rect 266360 33856 266412 33862
rect 266360 33798 266412 33804
rect 266268 18624 266320 18630
rect 266268 18566 266320 18572
rect 266372 3482 266400 33798
rect 266556 32570 266584 36910
rect 266544 32564 266596 32570
rect 266544 32506 266596 32512
rect 269040 21418 269068 43302
rect 270420 33794 270448 43302
rect 270500 40996 270552 41002
rect 270500 40938 270552 40944
rect 270408 33788 270460 33794
rect 270408 33730 270460 33736
rect 269028 21412 269080 21418
rect 269028 21354 269080 21360
rect 269120 19984 269172 19990
rect 269120 19926 269172 19932
rect 268108 3732 268160 3738
rect 268108 3674 268160 3680
rect 264992 3454 265848 3482
rect 266372 3454 267044 3482
rect 264612 3392 264664 3398
rect 264612 3334 264664 3340
rect 264624 480 264652 3334
rect 265820 480 265848 3454
rect 267016 480 267044 3454
rect 268120 480 268148 3674
rect 269132 3482 269160 19926
rect 269132 3454 269344 3482
rect 269316 480 269344 3454
rect 270512 3398 270540 40938
rect 271064 40118 271092 43316
rect 272260 41274 272288 43316
rect 272248 41268 272300 41274
rect 272248 41210 272300 41216
rect 273168 41268 273220 41274
rect 273168 41210 273220 41216
rect 271052 40112 271104 40118
rect 271052 40054 271104 40060
rect 272524 40112 272576 40118
rect 272524 40054 272576 40060
rect 272536 28354 272564 40054
rect 272524 28348 272576 28354
rect 272524 28290 272576 28296
rect 271880 24132 271932 24138
rect 271880 24074 271932 24080
rect 270592 6180 270644 6186
rect 270592 6122 270644 6128
rect 270500 3392 270552 3398
rect 270500 3334 270552 3340
rect 270604 3210 270632 6122
rect 271892 3482 271920 24074
rect 273180 19990 273208 41210
rect 273456 35358 273484 43316
rect 274652 40118 274680 43316
rect 275862 43302 275968 43330
rect 274640 40112 274692 40118
rect 274640 40054 274692 40060
rect 275836 40112 275888 40118
rect 275836 40054 275888 40060
rect 273260 35352 273312 35358
rect 273260 35294 273312 35300
rect 273444 35352 273496 35358
rect 273444 35294 273496 35300
rect 273168 19984 273220 19990
rect 273168 19926 273220 19932
rect 273272 3482 273300 35294
rect 275848 26994 275876 40054
rect 275836 26988 275888 26994
rect 275836 26930 275888 26936
rect 275940 24138 275968 43302
rect 277044 36650 277072 43316
rect 278254 43302 278728 43330
rect 279450 43302 280108 43330
rect 277032 36644 277084 36650
rect 277032 36586 277084 36592
rect 277400 36576 277452 36582
rect 277400 36518 277452 36524
rect 275928 24132 275980 24138
rect 275928 24074 275980 24080
rect 276020 22772 276072 22778
rect 276020 22714 276072 22720
rect 276032 3482 276060 22714
rect 271892 3454 272932 3482
rect 273272 3454 274128 3482
rect 276032 3454 276520 3482
rect 271696 3392 271748 3398
rect 271696 3334 271748 3340
rect 270512 3182 270632 3210
rect 270512 480 270540 3182
rect 271708 480 271736 3334
rect 272904 480 272932 3454
rect 274100 480 274128 3454
rect 275284 3324 275336 3330
rect 275284 3266 275336 3272
rect 275296 480 275324 3266
rect 276492 480 276520 3454
rect 277412 3380 277440 36518
rect 278700 22846 278728 43302
rect 278964 40724 279016 40730
rect 278964 40666 279016 40672
rect 278688 22840 278740 22846
rect 278688 22782 278740 22788
rect 278976 3482 279004 40666
rect 279976 6248 280028 6254
rect 279976 6190 280028 6196
rect 279988 6066 280016 6190
rect 280080 6186 280108 43302
rect 280632 38010 280660 43316
rect 281828 40118 281856 43316
rect 283024 40390 283052 43316
rect 284128 43302 284234 43330
rect 285430 43302 285628 43330
rect 286626 43302 287008 43330
rect 283012 40384 283064 40390
rect 283012 40326 283064 40332
rect 281816 40112 281868 40118
rect 281816 40054 281868 40060
rect 282828 40112 282880 40118
rect 282828 40054 282880 40060
rect 280160 38004 280212 38010
rect 280160 37946 280212 37952
rect 280620 38004 280672 38010
rect 280620 37946 280672 37952
rect 280068 6180 280120 6186
rect 280068 6122 280120 6128
rect 279988 6038 280108 6066
rect 278884 3454 279004 3482
rect 277412 3352 277716 3380
rect 277688 480 277716 3352
rect 278884 480 278912 3454
rect 280080 480 280108 6038
rect 280172 3380 280200 37946
rect 282840 6254 282868 40054
rect 284128 29646 284156 43302
rect 284208 40384 284260 40390
rect 284208 40326 284260 40332
rect 284116 29640 284168 29646
rect 284116 29582 284168 29588
rect 283656 7676 283708 7682
rect 283656 7618 283708 7624
rect 282828 6248 282880 6254
rect 282828 6190 282880 6196
rect 280172 3352 281304 3380
rect 281276 480 281304 3352
rect 282460 3120 282512 3126
rect 282460 3062 282512 3068
rect 282472 480 282500 3062
rect 283668 480 283696 7618
rect 284220 7614 284248 40326
rect 284300 29708 284352 29714
rect 284300 29650 284352 29656
rect 284208 7608 284260 7614
rect 284208 7550 284260 7556
rect 284312 3380 284340 29650
rect 285600 24206 285628 43302
rect 285772 40792 285824 40798
rect 285772 40734 285824 40740
rect 285588 24200 285640 24206
rect 285588 24142 285640 24148
rect 285784 3380 285812 40734
rect 286980 22778 287008 43302
rect 287808 39506 287836 43316
rect 289018 43302 289768 43330
rect 287796 39500 287848 39506
rect 287796 39442 287848 39448
rect 287060 39432 287112 39438
rect 287060 39374 287112 39380
rect 286968 22772 287020 22778
rect 286968 22714 287020 22720
rect 287072 3398 287100 39374
rect 287152 25560 287204 25566
rect 287152 25502 287204 25508
rect 287060 3392 287112 3398
rect 284312 3352 284800 3380
rect 285784 3352 285996 3380
rect 284772 480 284800 3352
rect 285968 480 285996 3352
rect 287060 3334 287112 3340
rect 287164 480 287192 25502
rect 289544 3936 289596 3942
rect 289544 3878 289596 3884
rect 288348 3392 288400 3398
rect 288348 3334 288400 3340
rect 288360 480 288388 3334
rect 289556 480 289584 3878
rect 289740 3806 289768 43302
rect 290200 40526 290228 43316
rect 290188 40520 290240 40526
rect 290188 40462 290240 40468
rect 291108 40520 291160 40526
rect 291108 40462 291160 40468
rect 291120 9042 291148 40462
rect 291396 40118 291424 43316
rect 292592 40118 292620 43316
rect 293710 43302 293816 43330
rect 294906 43302 295288 43330
rect 296102 43302 296668 43330
rect 297298 43302 298048 43330
rect 291384 40112 291436 40118
rect 291384 40054 291436 40060
rect 292488 40112 292540 40118
rect 292488 40054 292540 40060
rect 292580 40112 292632 40118
rect 292580 40054 292632 40060
rect 292500 31074 292528 40054
rect 291200 31068 291252 31074
rect 291200 31010 291252 31016
rect 292488 31068 292540 31074
rect 292488 31010 292540 31016
rect 290740 9036 290792 9042
rect 290740 8978 290792 8984
rect 291108 9036 291160 9042
rect 291108 8978 291160 8984
rect 289728 3800 289780 3806
rect 289728 3742 289780 3748
rect 290752 480 290780 8978
rect 291212 3482 291240 31010
rect 293788 25566 293816 43302
rect 293868 40112 293920 40118
rect 293868 40054 293920 40060
rect 293776 25560 293828 25566
rect 293776 25502 293828 25508
rect 293132 3596 293184 3602
rect 293132 3538 293184 3544
rect 291212 3454 291976 3482
rect 291948 480 291976 3454
rect 293144 480 293172 3538
rect 293880 3398 293908 40054
rect 295260 32502 295288 43302
rect 295248 32496 295300 32502
rect 295248 32438 295300 32444
rect 295340 32428 295392 32434
rect 295340 32370 295392 32376
rect 293960 10328 294012 10334
rect 293960 10270 294012 10276
rect 293972 3482 294000 10270
rect 295352 3482 295380 32370
rect 296640 3738 296668 43302
rect 296812 26920 296864 26926
rect 296812 26862 296864 26868
rect 296628 3732 296680 3738
rect 296628 3674 296680 3680
rect 296720 3664 296772 3670
rect 296720 3606 296772 3612
rect 293972 3454 294368 3482
rect 295352 3454 295564 3482
rect 293868 3392 293920 3398
rect 293868 3334 293920 3340
rect 294340 480 294368 3454
rect 295536 480 295564 3454
rect 296732 480 296760 3606
rect 296824 3210 296852 26862
rect 298020 10402 298048 43302
rect 298100 33924 298152 33930
rect 298100 33866 298152 33872
rect 298008 10396 298060 10402
rect 298008 10338 298060 10344
rect 298112 3210 298140 33866
rect 298480 33862 298508 43316
rect 299676 40594 299704 43316
rect 299664 40588 299716 40594
rect 299664 40530 299716 40536
rect 300768 40588 300820 40594
rect 300768 40530 300820 40536
rect 298468 33856 298520 33862
rect 298468 33798 298520 33804
rect 300308 4072 300360 4078
rect 300308 4014 300360 4020
rect 296824 3182 297956 3210
rect 298112 3182 299152 3210
rect 297928 480 297956 3182
rect 299124 480 299152 3182
rect 300320 480 300348 4014
rect 300780 3942 300808 40530
rect 300872 40526 300900 43316
rect 300860 40520 300912 40526
rect 300860 40462 300912 40468
rect 302068 35290 302096 43316
rect 303278 43302 303568 43330
rect 304474 43302 304948 43330
rect 302148 40520 302200 40526
rect 302148 40462 302200 40468
rect 302056 35284 302108 35290
rect 302056 35226 302108 35232
rect 302160 11762 302188 40462
rect 302240 35216 302292 35222
rect 302240 35158 302292 35164
rect 300860 11756 300912 11762
rect 300860 11698 300912 11704
rect 302148 11756 302200 11762
rect 302148 11698 302200 11704
rect 300768 3936 300820 3942
rect 300768 3878 300820 3884
rect 300872 2122 300900 11698
rect 302252 3210 302280 35158
rect 303540 4894 303568 43302
rect 304920 13122 304948 43302
rect 305656 36718 305684 43316
rect 306852 40118 306880 43316
rect 308048 40118 308076 43316
rect 309244 40118 309272 43316
rect 306840 40112 306892 40118
rect 306840 40054 306892 40060
rect 307668 40112 307720 40118
rect 307668 40054 307720 40060
rect 308036 40112 308088 40118
rect 308036 40054 308088 40060
rect 309048 40112 309100 40118
rect 309048 40054 309100 40060
rect 309232 40112 309284 40118
rect 309232 40054 309284 40060
rect 305000 36712 305052 36718
rect 305000 36654 305052 36660
rect 305644 36712 305696 36718
rect 305644 36654 305696 36660
rect 304908 13116 304960 13122
rect 304908 13058 304960 13064
rect 303528 4888 303580 4894
rect 303528 4830 303580 4836
rect 305012 3602 305040 36654
rect 305092 28280 305144 28286
rect 305092 28222 305144 28228
rect 305000 3596 305052 3602
rect 305000 3538 305052 3544
rect 305104 3482 305132 28222
rect 307392 4004 307444 4010
rect 307392 3946 307444 3952
rect 306196 3596 306248 3602
rect 306196 3538 306248 3544
rect 303804 3460 303856 3466
rect 303804 3402 303856 3408
rect 305012 3454 305132 3482
rect 302252 3182 302648 3210
rect 300872 2094 301452 2122
rect 301424 480 301452 2094
rect 302620 480 302648 3182
rect 303816 480 303844 3402
rect 305012 480 305040 3454
rect 306208 480 306236 3538
rect 307404 480 307432 3946
rect 307680 3466 307708 40054
rect 309060 14550 309088 40054
rect 309140 37936 309192 37942
rect 309140 37878 309192 37884
rect 309048 14544 309100 14550
rect 309048 14486 309100 14492
rect 307760 13184 307812 13190
rect 307760 13126 307812 13132
rect 307668 3460 307720 3466
rect 307668 3402 307720 3408
rect 307772 3346 307800 13126
rect 309152 3346 309180 37878
rect 310440 3602 310468 43316
rect 311650 43302 311848 43330
rect 311164 40112 311216 40118
rect 311164 40054 311216 40060
rect 311176 10470 311204 40054
rect 311820 26926 311848 43302
rect 312832 37942 312860 43316
rect 314042 43302 314608 43330
rect 313464 40384 313516 40390
rect 313464 40326 313516 40332
rect 312820 37936 312872 37942
rect 312820 37878 312872 37884
rect 311808 26920 311860 26926
rect 311808 26862 311860 26868
rect 311900 14476 311952 14482
rect 311900 14418 311952 14424
rect 311164 10464 311216 10470
rect 311164 10406 311216 10412
rect 310428 3596 310480 3602
rect 310428 3538 310480 3544
rect 310980 3528 311032 3534
rect 310980 3470 311032 3476
rect 307772 3318 308628 3346
rect 309152 3318 309824 3346
rect 308600 480 308628 3318
rect 309796 480 309824 3318
rect 310992 480 311020 3470
rect 311912 3346 311940 14418
rect 313372 4820 313424 4826
rect 313372 4762 313424 4768
rect 311912 3318 312216 3346
rect 312188 480 312216 3318
rect 313384 480 313412 4762
rect 313476 3346 313504 40326
rect 314580 3618 314608 43302
rect 315224 40118 315252 43316
rect 316420 40730 316448 43316
rect 316408 40724 316460 40730
rect 316408 40666 316460 40672
rect 317328 40724 317380 40730
rect 317328 40666 317380 40672
rect 315212 40112 315264 40118
rect 315212 40054 315264 40060
rect 315948 40112 316000 40118
rect 315948 40054 316000 40060
rect 315960 15978 315988 40054
rect 316040 29776 316092 29782
rect 316040 29718 316092 29724
rect 315948 15972 316000 15978
rect 315948 15914 316000 15920
rect 315764 4956 315816 4962
rect 315764 4898 315816 4904
rect 314580 3590 314700 3618
rect 313476 3318 314608 3346
rect 314580 480 314608 3318
rect 314672 3262 314700 3590
rect 314660 3256 314712 3262
rect 314660 3198 314712 3204
rect 315776 480 315804 4898
rect 316052 3346 316080 29718
rect 317340 25634 317368 40666
rect 317616 40118 317644 43316
rect 318720 41070 318748 43316
rect 318708 41064 318760 41070
rect 318708 41006 318760 41012
rect 317604 40112 317656 40118
rect 317604 40054 317656 40060
rect 318708 40112 318760 40118
rect 318708 40054 318760 40060
rect 317328 25628 317380 25634
rect 317328 25570 317380 25576
rect 318720 4010 318748 40054
rect 319916 39438 319944 43316
rect 321126 43302 321508 43330
rect 322322 43302 322888 43330
rect 319904 39432 319956 39438
rect 319904 39374 319956 39380
rect 320180 39364 320232 39370
rect 320180 39306 320232 39312
rect 318800 15904 318852 15910
rect 318800 15846 318852 15852
rect 318708 4004 318760 4010
rect 318708 3946 318760 3952
rect 318064 3868 318116 3874
rect 318064 3810 318116 3816
rect 316052 3318 317000 3346
rect 316972 480 317000 3318
rect 318076 480 318104 3810
rect 318812 3346 318840 15846
rect 320192 3346 320220 39306
rect 321480 3534 321508 43302
rect 321744 40860 321796 40866
rect 321744 40802 321796 40808
rect 321652 17264 321704 17270
rect 321652 17206 321704 17212
rect 321664 3670 321692 17206
rect 321652 3664 321704 3670
rect 321652 3606 321704 3612
rect 321468 3528 321520 3534
rect 321756 3482 321784 40802
rect 322860 17270 322888 43302
rect 323504 40118 323532 43316
rect 324700 40730 324728 43316
rect 324688 40724 324740 40730
rect 324688 40666 324740 40672
rect 325608 40724 325660 40730
rect 325608 40666 325660 40672
rect 323492 40112 323544 40118
rect 323492 40054 323544 40060
rect 324228 40112 324280 40118
rect 324228 40054 324280 40060
rect 324240 31142 324268 40054
rect 322940 31136 322992 31142
rect 322940 31078 322992 31084
rect 324228 31136 324280 31142
rect 324228 31078 324280 31084
rect 322848 17264 322900 17270
rect 322848 17206 322900 17212
rect 322848 3664 322900 3670
rect 322848 3606 322900 3612
rect 321468 3470 321520 3476
rect 321664 3454 321784 3482
rect 318812 3318 319300 3346
rect 320192 3318 320496 3346
rect 319272 480 319300 3318
rect 320468 480 320496 3318
rect 321664 480 321692 3454
rect 322860 480 322888 3606
rect 322952 3346 322980 31078
rect 325240 4140 325292 4146
rect 325240 4082 325292 4088
rect 322952 3318 324084 3346
rect 324056 480 324084 3318
rect 325252 480 325280 4082
rect 325620 3874 325648 40666
rect 325896 40118 325924 43316
rect 325884 40112 325936 40118
rect 325884 40054 325936 40060
rect 326988 40112 327040 40118
rect 326988 40054 327040 40060
rect 327000 18630 327028 40054
rect 327092 36938 327120 43316
rect 328302 43302 328408 43330
rect 329498 43302 329788 43330
rect 330694 43302 331168 43330
rect 331890 43302 332548 43330
rect 327092 36910 327304 36938
rect 327080 32564 327132 32570
rect 327080 32506 327132 32512
rect 325700 18624 325752 18630
rect 325700 18566 325752 18572
rect 326988 18624 327040 18630
rect 326988 18566 327040 18572
rect 325608 3868 325660 3874
rect 325608 3810 325660 3816
rect 325712 3346 325740 18566
rect 327092 3346 327120 32506
rect 327276 32434 327304 36910
rect 327264 32428 327316 32434
rect 327264 32370 327316 32376
rect 328380 3670 328408 43302
rect 328552 40928 328604 40934
rect 328552 40870 328604 40876
rect 328368 3664 328420 3670
rect 328368 3606 328420 3612
rect 328564 3346 328592 40870
rect 329760 28286 329788 43302
rect 329748 28280 329800 28286
rect 329748 28222 329800 28228
rect 329840 21412 329892 21418
rect 329840 21354 329892 21360
rect 329852 3346 329880 21354
rect 331140 11830 331168 43302
rect 331220 33788 331272 33794
rect 331220 33730 331272 33736
rect 331128 11824 331180 11830
rect 331128 11766 331180 11772
rect 325712 3318 326476 3346
rect 327092 3318 327672 3346
rect 328564 3318 328868 3346
rect 329852 3318 330064 3346
rect 326448 480 326476 3318
rect 327644 480 327672 3318
rect 328840 480 328868 3318
rect 330036 480 330064 3318
rect 331232 480 331260 33730
rect 331312 28348 331364 28354
rect 331312 28290 331364 28296
rect 331324 3346 331352 28290
rect 331324 3318 332456 3346
rect 332428 480 332456 3318
rect 332520 3194 332548 43302
rect 333072 40798 333100 43316
rect 334268 40798 334296 43316
rect 333060 40792 333112 40798
rect 333060 40734 333112 40740
rect 333888 40792 333940 40798
rect 333888 40734 333940 40740
rect 334256 40792 334308 40798
rect 334256 40734 334308 40740
rect 333900 19990 333928 40734
rect 335464 40390 335492 43316
rect 336568 43302 336674 43330
rect 337870 43302 338068 43330
rect 339066 43302 339448 43330
rect 340262 43302 340828 43330
rect 341458 43302 342208 43330
rect 335452 40384 335504 40390
rect 335452 40326 335504 40332
rect 333980 35352 334032 35358
rect 333980 35294 334032 35300
rect 332600 19984 332652 19990
rect 332600 19926 332652 19932
rect 333888 19984 333940 19990
rect 333888 19926 333940 19932
rect 332612 3346 332640 19926
rect 333992 3346 334020 35294
rect 335360 26988 335412 26994
rect 335360 26930 335412 26936
rect 335372 3482 335400 26930
rect 336568 21418 336596 43302
rect 336648 40384 336700 40390
rect 336648 40326 336700 40332
rect 336556 21412 336608 21418
rect 336556 21354 336608 21360
rect 335372 3454 335952 3482
rect 332612 3318 333652 3346
rect 333992 3318 334756 3346
rect 332508 3188 332560 3194
rect 332508 3130 332560 3136
rect 333624 480 333652 3318
rect 334728 480 334756 3318
rect 335924 480 335952 3454
rect 336660 3126 336688 40326
rect 338040 33794 338068 43302
rect 338120 36644 338172 36650
rect 338120 36586 338172 36592
rect 338028 33788 338080 33794
rect 338028 33730 338080 33736
rect 336740 24132 336792 24138
rect 336740 24074 336792 24080
rect 336752 3482 336780 24074
rect 338132 3482 338160 36586
rect 336752 3454 337148 3482
rect 338132 3454 338344 3482
rect 336648 3120 336700 3126
rect 336648 3062 336700 3068
rect 337120 480 337148 3454
rect 338316 480 338344 3454
rect 339420 3369 339448 43302
rect 339500 22840 339552 22846
rect 339500 22782 339552 22788
rect 339406 3360 339462 3369
rect 339406 3295 339462 3304
rect 339512 480 339540 22782
rect 340800 7682 340828 43302
rect 340880 38004 340932 38010
rect 340880 37946 340932 37952
rect 340788 7676 340840 7682
rect 340788 7618 340840 7624
rect 340696 6180 340748 6186
rect 340696 6122 340748 6128
rect 340708 480 340736 6122
rect 340892 3482 340920 37946
rect 342180 35222 342208 43302
rect 342640 40118 342668 43316
rect 343744 41070 343772 43316
rect 343732 41064 343784 41070
rect 343732 41006 343784 41012
rect 344836 41064 344888 41070
rect 344836 41006 344888 41012
rect 342628 40112 342680 40118
rect 342628 40054 342680 40060
rect 343548 40112 343600 40118
rect 343548 40054 343600 40060
rect 342168 35216 342220 35222
rect 342168 35158 342220 35164
rect 343088 6248 343140 6254
rect 343088 6190 343140 6196
rect 340892 3454 341932 3482
rect 341904 480 341932 3454
rect 343100 480 343128 6190
rect 343560 3330 343588 40054
rect 344848 24138 344876 41006
rect 344836 24132 344888 24138
rect 344836 24074 344888 24080
rect 344940 14482 344968 43316
rect 345664 40928 345716 40934
rect 345664 40870 345716 40876
rect 345020 29640 345072 29646
rect 345020 29582 345072 29588
rect 344928 14476 344980 14482
rect 344928 14418 344980 14424
rect 344284 7608 344336 7614
rect 344284 7550 344336 7556
rect 343548 3324 343600 3330
rect 343548 3266 343600 3272
rect 344296 480 344324 7550
rect 345032 3482 345060 29582
rect 345676 6186 345704 40870
rect 346136 40730 346164 43316
rect 347346 43302 347728 43330
rect 346124 40724 346176 40730
rect 346124 40666 346176 40672
rect 346400 24200 346452 24206
rect 346400 24142 346452 24148
rect 345664 6180 345716 6186
rect 345664 6122 345716 6128
rect 346412 3482 346440 24142
rect 347700 8974 347728 43302
rect 347780 39500 347832 39506
rect 347780 39442 347832 39448
rect 347688 8968 347740 8974
rect 347688 8910 347740 8916
rect 345032 3454 345520 3482
rect 346412 3454 346716 3482
rect 345492 480 345520 3454
rect 346688 480 346716 3454
rect 347792 2106 347820 39442
rect 348528 36582 348556 43316
rect 349738 43302 350488 43330
rect 348516 36576 348568 36582
rect 348516 36518 348568 36524
rect 347872 22772 347924 22778
rect 347872 22714 347924 22720
rect 347780 2100 347832 2106
rect 347780 2042 347832 2048
rect 347884 480 347912 22714
rect 350460 4078 350488 43302
rect 350920 40118 350948 43316
rect 352116 40118 352144 43316
rect 353312 40118 353340 43316
rect 350908 40112 350960 40118
rect 350908 40054 350960 40060
rect 351828 40112 351880 40118
rect 351828 40054 351880 40060
rect 352104 40112 352156 40118
rect 352104 40054 352156 40060
rect 353208 40112 353260 40118
rect 353208 40054 353260 40060
rect 353300 40112 353352 40118
rect 353300 40054 353352 40060
rect 351840 22778 351868 40054
rect 351920 31068 351972 31074
rect 351920 31010 351972 31016
rect 351828 22772 351880 22778
rect 351828 22714 351880 22720
rect 351368 9036 351420 9042
rect 351368 8978 351420 8984
rect 350448 4072 350500 4078
rect 350448 4014 350500 4020
rect 350264 3800 350316 3806
rect 350264 3742 350316 3748
rect 349068 2100 349120 2106
rect 349068 2042 349120 2048
rect 349080 480 349108 2042
rect 350276 480 350304 3742
rect 351380 480 351408 8978
rect 351932 3482 351960 31010
rect 353220 26994 353248 40054
rect 354508 29646 354536 43316
rect 355718 43302 356008 43330
rect 356914 43302 357388 43330
rect 358110 43302 358768 43330
rect 354588 40112 354640 40118
rect 354588 40054 354640 40060
rect 354496 29640 354548 29646
rect 354496 29582 354548 29588
rect 353208 26988 353260 26994
rect 353208 26930 353260 26936
rect 354600 3806 354628 40054
rect 354680 25560 354732 25566
rect 354680 25502 354732 25508
rect 354588 3800 354640 3806
rect 354588 3742 354640 3748
rect 351932 3454 352604 3482
rect 352576 480 352604 3454
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 354692 3346 354720 25502
rect 355980 10334 356008 43302
rect 356152 32496 356204 32502
rect 356152 32438 356204 32444
rect 355968 10328 356020 10334
rect 355968 10270 356020 10276
rect 353772 480 353800 3334
rect 354692 3318 354996 3346
rect 354968 480 354996 3318
rect 356164 480 356192 32438
rect 357360 5114 357388 43302
rect 357440 10396 357492 10402
rect 357440 10338 357492 10344
rect 357176 5086 357388 5114
rect 357176 3398 357204 5086
rect 357348 3732 357400 3738
rect 357348 3674 357400 3680
rect 357164 3392 357216 3398
rect 357164 3334 357216 3340
rect 357360 480 357388 3674
rect 357452 3346 357480 10338
rect 358740 5166 358768 43302
rect 359292 38010 359320 43316
rect 360488 40118 360516 43316
rect 361684 40118 361712 43316
rect 362788 43302 362894 43330
rect 364090 43302 364288 43330
rect 365286 43302 365668 43330
rect 360476 40112 360528 40118
rect 360476 40054 360528 40060
rect 361488 40112 361540 40118
rect 361488 40054 361540 40060
rect 361672 40112 361724 40118
rect 361672 40054 361724 40060
rect 359280 38004 359332 38010
rect 359280 37946 359332 37952
rect 358820 33856 358872 33862
rect 358820 33798 358872 33804
rect 358728 5160 358780 5166
rect 358728 5102 358780 5108
rect 358832 3346 358860 33798
rect 360936 3936 360988 3942
rect 360936 3878 360988 3884
rect 357452 3318 358584 3346
rect 358832 3318 359780 3346
rect 358556 480 358584 3318
rect 359752 480 359780 3318
rect 360948 480 360976 3878
rect 361500 3738 361528 40054
rect 362788 25566 362816 43302
rect 362868 40112 362920 40118
rect 362868 40054 362920 40060
rect 362776 25560 362828 25566
rect 362776 25502 362828 25508
rect 361580 11756 361632 11762
rect 361580 11698 361632 11704
rect 361488 3732 361540 3738
rect 361488 3674 361540 3680
rect 361592 1986 361620 11698
rect 362880 5030 362908 40054
rect 362960 35284 363012 35290
rect 362960 35226 363012 35232
rect 362868 5024 362920 5030
rect 362868 4966 362920 4972
rect 362972 3346 363000 35226
rect 364260 3505 364288 43302
rect 365640 5370 365668 43302
rect 366468 39370 366496 43316
rect 367664 41070 367692 43316
rect 367652 41064 367704 41070
rect 367652 41006 367704 41012
rect 367744 40792 367796 40798
rect 367744 40734 367796 40740
rect 366456 39364 366508 39370
rect 366456 39306 366508 39312
rect 365720 36712 365772 36718
rect 365720 36654 365772 36660
rect 365628 5364 365680 5370
rect 365628 5306 365680 5312
rect 364524 4888 364576 4894
rect 364524 4830 364576 4836
rect 364246 3496 364302 3505
rect 364246 3431 364302 3440
rect 362972 3318 363368 3346
rect 361592 1958 362172 1986
rect 362144 480 362172 1958
rect 363340 480 363368 3318
rect 364536 480 364564 4830
rect 365732 3466 365760 36654
rect 367756 13190 367784 40734
rect 368860 40118 368888 43316
rect 369964 41274 369992 43316
rect 369952 41268 370004 41274
rect 369952 41210 370004 41216
rect 371056 41268 371108 41274
rect 371056 41210 371108 41216
rect 368848 40112 368900 40118
rect 368848 40054 368900 40060
rect 369768 40112 369820 40118
rect 369768 40054 369820 40060
rect 368480 14544 368532 14550
rect 368480 14486 368532 14492
rect 367744 13184 367796 13190
rect 367744 13126 367796 13132
rect 365812 13116 365864 13122
rect 365812 13058 365864 13064
rect 365720 3460 365772 3466
rect 365720 3402 365772 3408
rect 365824 1442 365852 13058
rect 368020 3596 368072 3602
rect 368020 3538 368072 3544
rect 366916 3460 366968 3466
rect 366916 3402 366968 3408
rect 365732 1414 365852 1442
rect 365732 480 365760 1414
rect 366928 480 366956 3402
rect 368032 480 368060 3538
rect 368492 3346 368520 14486
rect 369780 5438 369808 40054
rect 371068 31074 371096 41210
rect 371056 31068 371108 31074
rect 371056 31010 371108 31016
rect 370412 10464 370464 10470
rect 370412 10406 370464 10412
rect 369768 5432 369820 5438
rect 369768 5374 369820 5380
rect 368492 3318 369256 3346
rect 369228 480 369256 3318
rect 370424 480 370452 10406
rect 371160 3466 371188 43316
rect 372370 43302 372568 43330
rect 373566 43302 373948 43330
rect 372540 4826 372568 43302
rect 373920 32502 373948 43302
rect 374748 40934 374776 43316
rect 374736 40928 374788 40934
rect 374736 40870 374788 40876
rect 375944 40118 375972 43316
rect 377140 40118 377168 43316
rect 378336 40662 378364 43316
rect 378324 40656 378376 40662
rect 378324 40598 378376 40604
rect 379428 40656 379480 40662
rect 379428 40598 379480 40604
rect 375932 40112 375984 40118
rect 375932 40054 375984 40060
rect 376668 40112 376720 40118
rect 376668 40054 376720 40060
rect 377128 40112 377180 40118
rect 377128 40054 377180 40060
rect 378048 40112 378100 40118
rect 378048 40054 378100 40060
rect 374092 37936 374144 37942
rect 374092 37878 374144 37884
rect 373908 32496 373960 32502
rect 373908 32438 373960 32444
rect 372712 26920 372764 26926
rect 372712 26862 372764 26868
rect 372724 19394 372752 26862
rect 372632 19366 372752 19394
rect 372632 19310 372660 19366
rect 372620 19304 372672 19310
rect 372620 19246 372672 19252
rect 372804 12300 372856 12306
rect 372804 12242 372856 12248
rect 372528 4820 372580 4826
rect 372528 4762 372580 4768
rect 371148 3460 371200 3466
rect 371148 3402 371200 3408
rect 371608 3052 371660 3058
rect 371608 2994 371660 3000
rect 371620 480 371648 2994
rect 372816 480 372844 12242
rect 374104 592 374132 37878
rect 375380 15972 375432 15978
rect 375380 15914 375432 15920
rect 375196 3256 375248 3262
rect 375196 3198 375248 3204
rect 374012 564 374132 592
rect 374012 480 374040 564
rect 375208 480 375236 3198
rect 375392 610 375420 15914
rect 376680 5234 376708 40054
rect 378060 28354 378088 40054
rect 378048 28348 378100 28354
rect 378048 28290 378100 28296
rect 376760 25628 376812 25634
rect 376760 25570 376812 25576
rect 376668 5228 376720 5234
rect 376668 5170 376720 5176
rect 376772 610 376800 25570
rect 379440 4146 379468 40598
rect 379532 40118 379560 43316
rect 379520 40112 379572 40118
rect 379520 40054 379572 40060
rect 380728 11762 380756 43316
rect 381924 40866 381952 43316
rect 383488 41426 383516 43438
rect 384330 43302 384988 43330
rect 383488 41398 383608 41426
rect 381912 40860 381964 40866
rect 381912 40802 381964 40808
rect 380808 40112 380860 40118
rect 380808 40054 380860 40060
rect 380716 11756 380768 11762
rect 380716 11698 380768 11704
rect 379980 6180 380032 6186
rect 379980 6122 380032 6128
rect 379428 4140 379480 4146
rect 379428 4082 379480 4088
rect 378784 4004 378836 4010
rect 378784 3946 378836 3952
rect 375380 604 375432 610
rect 375380 546 375432 552
rect 376392 604 376444 610
rect 376392 546 376444 552
rect 376760 604 376812 610
rect 376760 546 376812 552
rect 377588 604 377640 610
rect 377588 546 377640 552
rect 376404 480 376432 546
rect 377600 480 377628 546
rect 378796 480 378824 3946
rect 379992 480 380020 6122
rect 380820 5506 380848 40054
rect 380900 39432 380952 39438
rect 380900 39374 380952 39380
rect 380808 5500 380860 5506
rect 380808 5442 380860 5448
rect 380912 626 380940 39374
rect 383580 33862 383608 41398
rect 384960 33862 384988 43302
rect 385512 40118 385540 43316
rect 386708 40118 386736 43316
rect 387904 40118 387932 43316
rect 389100 40798 389128 43316
rect 390310 43302 390508 43330
rect 391506 43302 391888 43330
rect 392702 43302 393268 43330
rect 393898 43302 394648 43330
rect 389088 40792 389140 40798
rect 389088 40734 389140 40740
rect 385500 40112 385552 40118
rect 385500 40054 385552 40060
rect 386328 40112 386380 40118
rect 386328 40054 386380 40060
rect 386696 40112 386748 40118
rect 386696 40054 386748 40060
rect 387708 40112 387760 40118
rect 387708 40054 387760 40060
rect 387892 40112 387944 40118
rect 387892 40054 387944 40060
rect 389088 40112 389140 40118
rect 389088 40054 389140 40060
rect 383108 33856 383160 33862
rect 383108 33798 383160 33804
rect 383568 33856 383620 33862
rect 383568 33798 383620 33804
rect 384948 33856 385000 33862
rect 384948 33798 385000 33804
rect 383120 29073 383148 33798
rect 383660 31136 383712 31142
rect 383660 31078 383712 31084
rect 383106 29064 383162 29073
rect 383106 28999 383162 29008
rect 383290 29064 383346 29073
rect 383290 28999 383346 29008
rect 383304 28966 383332 28999
rect 383292 28960 383344 28966
rect 383292 28902 383344 28908
rect 383476 22024 383528 22030
rect 383476 21966 383528 21972
rect 382372 17264 382424 17270
rect 382372 17206 382424 17212
rect 382384 7614 382412 17206
rect 383488 12442 383516 21966
rect 383292 12436 383344 12442
rect 383292 12378 383344 12384
rect 383476 12436 383528 12442
rect 383476 12378 383528 12384
rect 382372 7608 382424 7614
rect 382372 7550 382424 7556
rect 383304 4962 383332 12378
rect 383568 7608 383620 7614
rect 383568 7550 383620 7556
rect 383292 4956 383344 4962
rect 383292 4898 383344 4904
rect 382372 3528 382424 3534
rect 382372 3470 382424 3476
rect 380912 598 381124 626
rect 381096 592 381124 598
rect 381096 564 381216 592
rect 381188 480 381216 564
rect 382384 480 382412 3470
rect 383580 480 383608 7550
rect 383672 610 383700 31078
rect 386340 4010 386368 40054
rect 386420 18624 386472 18630
rect 386420 18566 386472 18572
rect 386328 4004 386380 4010
rect 386328 3946 386380 3952
rect 385868 3868 385920 3874
rect 385868 3810 385920 3816
rect 383660 604 383712 610
rect 383660 546 383712 552
rect 384672 604 384724 610
rect 384672 546 384724 552
rect 384684 480 384712 546
rect 385880 480 385908 3810
rect 386432 610 386460 18566
rect 387720 5302 387748 40054
rect 387800 32428 387852 32434
rect 387800 32370 387852 32376
rect 387708 5296 387760 5302
rect 387708 5238 387760 5244
rect 387812 610 387840 32370
rect 389100 13122 389128 40054
rect 390376 19304 390428 19310
rect 390376 19246 390428 19252
rect 389088 13116 389140 13122
rect 389088 13058 389140 13064
rect 390388 9761 390416 19246
rect 390374 9752 390430 9761
rect 390374 9687 390430 9696
rect 390480 4894 390508 43302
rect 391860 35290 391888 43302
rect 391848 35284 391900 35290
rect 391848 35226 391900 35232
rect 390560 28280 390612 28286
rect 390560 28222 390612 28228
rect 390572 19310 390600 28222
rect 390560 19304 390612 19310
rect 390560 19246 390612 19252
rect 391848 11824 391900 11830
rect 391848 11766 391900 11772
rect 390650 9752 390706 9761
rect 390650 9687 390706 9696
rect 390664 9654 390692 9687
rect 390652 9648 390704 9654
rect 390652 9590 390704 9596
rect 390652 9512 390704 9518
rect 390652 9454 390704 9460
rect 390468 4888 390520 4894
rect 390468 4830 390520 4836
rect 389456 3664 389508 3670
rect 389456 3606 389508 3612
rect 386420 604 386472 610
rect 386420 546 386472 552
rect 387064 604 387116 610
rect 387064 546 387116 552
rect 387800 604 387852 610
rect 387800 546 387852 552
rect 388260 604 388312 610
rect 388260 546 388312 552
rect 387076 480 387104 546
rect 388272 480 388300 546
rect 389468 480 389496 3606
rect 390664 480 390692 9454
rect 391860 480 391888 11766
rect 393240 3942 393268 43302
rect 393320 19984 393372 19990
rect 393320 19926 393372 19932
rect 393228 3936 393280 3942
rect 393228 3878 393280 3884
rect 393044 3188 393096 3194
rect 393044 3130 393096 3136
rect 393056 480 393084 3130
rect 393332 2854 393360 19926
rect 394620 5098 394648 43302
rect 394988 40118 395016 43316
rect 396184 41138 396212 43316
rect 396172 41132 396224 41138
rect 396172 41074 396224 41080
rect 394976 40112 395028 40118
rect 394976 40054 395028 40060
rect 395988 40112 396040 40118
rect 395988 40054 396040 40060
rect 396000 14550 396028 40054
rect 397380 15910 397408 43316
rect 398590 43302 398788 43330
rect 399786 43302 400168 43330
rect 400982 43302 401548 43330
rect 397460 21412 397512 21418
rect 397460 21354 397512 21360
rect 397368 15904 397420 15910
rect 397368 15846 397420 15852
rect 395988 14544 396040 14550
rect 395988 14486 396040 14492
rect 394700 13184 394752 13190
rect 394700 13126 394752 13132
rect 394608 5092 394660 5098
rect 394608 5034 394660 5040
rect 394712 2854 394740 13126
rect 396632 3120 396684 3126
rect 396632 3062 396684 3068
rect 393320 2848 393372 2854
rect 393320 2790 393372 2796
rect 394700 2848 394752 2854
rect 394700 2790 394752 2796
rect 394240 2780 394292 2786
rect 394240 2722 394292 2728
rect 395436 2780 395488 2786
rect 395436 2722 395488 2728
rect 394252 480 394280 2722
rect 395448 480 395476 2722
rect 396644 480 396672 3062
rect 397472 2854 397500 21354
rect 398760 6186 398788 43302
rect 398932 33788 398984 33794
rect 398932 33730 398984 33736
rect 398944 29050 398972 33730
rect 398852 29022 398972 29050
rect 398852 27606 398880 29022
rect 398840 27600 398892 27606
rect 398840 27542 398892 27548
rect 398932 27600 398984 27606
rect 398932 27542 398984 27548
rect 398748 6180 398800 6186
rect 398748 6122 398800 6128
rect 398944 4842 398972 27542
rect 398944 4814 399064 4842
rect 397460 2848 397512 2854
rect 397460 2790 397512 2796
rect 397828 2780 397880 2786
rect 397828 2722 397880 2728
rect 397840 480 397868 2722
rect 399036 480 399064 4814
rect 400140 3874 400168 43302
rect 401520 17338 401548 43302
rect 402164 38078 402192 43316
rect 403360 41070 403388 43316
rect 403348 41064 403400 41070
rect 403348 41006 403400 41012
rect 404556 40118 404584 43316
rect 405752 40118 405780 43316
rect 406962 43302 407068 43330
rect 408158 43302 408448 43330
rect 409354 43302 409828 43330
rect 410550 43302 411208 43330
rect 404544 40112 404596 40118
rect 404544 40054 404596 40060
rect 405648 40112 405700 40118
rect 405648 40054 405700 40060
rect 405740 40112 405792 40118
rect 405740 40054 405792 40060
rect 406936 40112 406988 40118
rect 406936 40054 406988 40060
rect 402152 38072 402204 38078
rect 402152 38014 402204 38020
rect 401600 35216 401652 35222
rect 401600 35158 401652 35164
rect 401508 17332 401560 17338
rect 401508 17274 401560 17280
rect 401612 12442 401640 35158
rect 404360 24132 404412 24138
rect 404360 24074 404412 24080
rect 404372 12442 404400 24074
rect 405660 19990 405688 40054
rect 406948 29714 406976 40054
rect 406936 29708 406988 29714
rect 406936 29650 406988 29656
rect 405648 19984 405700 19990
rect 405648 19926 405700 19932
rect 405740 14476 405792 14482
rect 405740 14418 405792 14424
rect 401600 12436 401652 12442
rect 401600 12378 401652 12384
rect 402520 12436 402572 12442
rect 402520 12378 402572 12384
rect 404360 12436 404412 12442
rect 404360 12378 404412 12384
rect 404912 12436 404964 12442
rect 404912 12378 404964 12384
rect 401324 7676 401376 7682
rect 401324 7618 401376 7624
rect 400128 3868 400180 3874
rect 400128 3810 400180 3816
rect 400218 3360 400274 3369
rect 400218 3295 400274 3304
rect 400232 480 400260 3295
rect 401336 480 401364 7618
rect 402532 480 402560 12378
rect 403716 3324 403768 3330
rect 403716 3266 403768 3272
rect 403728 480 403756 3266
rect 404924 480 404952 12378
rect 405752 610 405780 14418
rect 407040 3369 407068 43302
rect 407212 40724 407264 40730
rect 407212 40666 407264 40672
rect 407026 3360 407082 3369
rect 407026 3295 407082 3304
rect 407224 626 407252 40666
rect 408420 18630 408448 43302
rect 408500 36576 408552 36582
rect 408500 36518 408552 36524
rect 408408 18624 408460 18630
rect 408408 18566 408460 18572
rect 408512 7614 408540 36518
rect 409800 26926 409828 43302
rect 409788 26920 409840 26926
rect 409788 26862 409840 26868
rect 408592 8968 408644 8974
rect 408592 8910 408644 8916
rect 408500 7608 408552 7614
rect 408500 7550 408552 7556
rect 408604 7426 408632 8910
rect 409696 7608 409748 7614
rect 409696 7550 409748 7556
rect 408512 7398 408632 7426
rect 405740 604 405792 610
rect 405740 546 405792 552
rect 406108 604 406160 610
rect 407224 598 407344 626
rect 406108 546 406160 552
rect 406120 480 406148 546
rect 407316 480 407344 598
rect 408512 480 408540 7398
rect 409708 480 409736 7550
rect 411180 4078 411208 43302
rect 411732 40118 411760 43316
rect 412928 40118 412956 43316
rect 414124 40118 414152 43316
rect 415228 43302 415334 43330
rect 416530 43302 416728 43330
rect 417726 43302 418108 43330
rect 418922 43302 419488 43330
rect 411720 40112 411772 40118
rect 411720 40054 411772 40060
rect 412548 40112 412600 40118
rect 412548 40054 412600 40060
rect 412916 40112 412968 40118
rect 412916 40054 412968 40060
rect 413928 40112 413980 40118
rect 413928 40054 413980 40060
rect 414112 40112 414164 40118
rect 414112 40054 414164 40060
rect 412560 22778 412588 40054
rect 413940 35222 413968 40054
rect 415228 36582 415256 43302
rect 415308 40112 415360 40118
rect 415308 40054 415360 40060
rect 415216 36576 415268 36582
rect 415216 36518 415268 36524
rect 413928 35216 413980 35222
rect 413928 35158 413980 35164
rect 411260 22772 411312 22778
rect 411260 22714 411312 22720
rect 412548 22772 412600 22778
rect 412548 22714 412600 22720
rect 411272 9654 411300 22714
rect 412640 19372 412692 19378
rect 412640 19314 412692 19320
rect 411260 9648 411312 9654
rect 411260 9590 411312 9596
rect 410892 4072 410944 4078
rect 410892 4014 410944 4020
rect 411168 4072 411220 4078
rect 411168 4014 411220 4020
rect 410904 480 410932 4014
rect 412652 2854 412680 19314
rect 414480 3800 414532 3806
rect 414480 3742 414532 3748
rect 412640 2848 412692 2854
rect 412640 2790 412692 2796
rect 413284 2780 413336 2786
rect 413284 2722 413336 2728
rect 412088 604 412140 610
rect 412088 546 412140 552
rect 412100 480 412128 546
rect 413296 480 413324 2722
rect 414492 480 414520 3742
rect 415320 3602 415348 40054
rect 415400 29640 415452 29646
rect 415400 29582 415452 29588
rect 415412 9654 415440 29582
rect 416700 10402 416728 43302
rect 416688 10396 416740 10402
rect 416688 10338 416740 10344
rect 416872 10328 416924 10334
rect 416872 10270 416924 10276
rect 415400 9648 415452 9654
rect 415400 9590 415452 9596
rect 415308 3596 415360 3602
rect 415308 3538 415360 3544
rect 415676 604 415728 610
rect 415676 546 415728 552
rect 415688 480 415716 546
rect 416884 480 416912 10270
rect 418080 3670 418108 43302
rect 419460 21486 419488 43302
rect 420104 40118 420132 43316
rect 421208 40118 421236 43316
rect 422404 40118 422432 43316
rect 423508 43302 423614 43330
rect 424810 43302 425008 43330
rect 426006 43302 426388 43330
rect 427202 43302 427768 43330
rect 420092 40112 420144 40118
rect 420092 40054 420144 40060
rect 420828 40112 420880 40118
rect 420828 40054 420880 40060
rect 421196 40112 421248 40118
rect 421196 40054 421248 40060
rect 422208 40112 422260 40118
rect 422208 40054 422260 40060
rect 422392 40112 422444 40118
rect 422392 40054 422444 40060
rect 419540 38004 419592 38010
rect 419540 37946 419592 37952
rect 419448 21480 419500 21486
rect 419448 21422 419500 21428
rect 419172 5160 419224 5166
rect 419172 5102 419224 5108
rect 418068 3664 418120 3670
rect 418068 3606 418120 3612
rect 417976 3392 418028 3398
rect 417976 3334 418028 3340
rect 417988 480 418016 3334
rect 419184 480 419212 5102
rect 419552 2854 419580 37946
rect 420840 32434 420868 40054
rect 420828 32428 420880 32434
rect 420828 32370 420880 32376
rect 422220 3738 422248 40054
rect 423508 24138 423536 43302
rect 423588 40112 423640 40118
rect 423588 40054 423640 40060
rect 423496 24132 423548 24138
rect 423496 24074 423548 24080
rect 423600 6254 423628 40054
rect 423680 25560 423732 25566
rect 423680 25502 423732 25508
rect 423588 6248 423640 6254
rect 423588 6190 423640 6196
rect 422760 5024 422812 5030
rect 422760 4966 422812 4972
rect 421564 3732 421616 3738
rect 421564 3674 421616 3680
rect 422208 3732 422260 3738
rect 422208 3674 422260 3680
rect 419540 2848 419592 2854
rect 419540 2790 419592 2796
rect 420368 2780 420420 2786
rect 420368 2722 420420 2728
rect 420380 480 420408 2722
rect 421576 480 421604 3674
rect 422772 480 422800 4966
rect 423692 2802 423720 25502
rect 424980 15978 425008 43302
rect 424968 15972 425020 15978
rect 424968 15914 425020 15920
rect 426360 7614 426388 43302
rect 426440 39364 426492 39370
rect 426440 39306 426492 39312
rect 426348 7608 426400 7614
rect 426348 7550 426400 7556
rect 426348 5364 426400 5370
rect 426348 5306 426400 5312
rect 425058 4856 425114 4865
rect 425058 4791 425060 4800
rect 425112 4791 425114 4800
rect 425060 4762 425112 4768
rect 425150 3496 425206 3505
rect 425150 3431 425206 3440
rect 423692 2774 423904 2802
rect 423876 2666 423904 2774
rect 423876 2638 423996 2666
rect 423968 480 423996 2638
rect 425164 480 425192 3431
rect 426360 480 426388 5306
rect 426452 2854 426480 39306
rect 427740 25634 427768 43302
rect 427912 40996 427964 41002
rect 427912 40938 427964 40944
rect 427728 25628 427780 25634
rect 427728 25570 427780 25576
rect 427924 2854 427952 40938
rect 428384 40118 428412 43316
rect 429580 40118 429608 43316
rect 430776 40118 430804 43316
rect 431972 40118 432000 43316
rect 433182 43302 433288 43330
rect 434378 43302 434668 43330
rect 435574 43302 436048 43330
rect 436770 43302 437428 43330
rect 428372 40112 428424 40118
rect 428372 40054 428424 40060
rect 429108 40112 429160 40118
rect 429108 40054 429160 40060
rect 429568 40112 429620 40118
rect 429568 40054 429620 40060
rect 430488 40112 430540 40118
rect 430488 40054 430540 40060
rect 430764 40112 430816 40118
rect 430764 40054 430816 40060
rect 431868 40112 431920 40118
rect 431868 40054 431920 40060
rect 431960 40112 432012 40118
rect 431960 40054 432012 40060
rect 433156 40112 433208 40118
rect 433156 40054 433208 40060
rect 429120 3534 429148 40054
rect 430500 8974 430528 40054
rect 430580 31068 430632 31074
rect 430580 31010 430632 31016
rect 430488 8968 430540 8974
rect 430488 8910 430540 8916
rect 429936 5432 429988 5438
rect 429936 5374 429988 5380
rect 429108 3528 429160 3534
rect 429108 3470 429160 3476
rect 426440 2848 426492 2854
rect 426440 2790 426492 2796
rect 427912 2848 427964 2854
rect 427912 2790 427964 2796
rect 427544 2780 427596 2786
rect 427544 2722 427596 2728
rect 428740 2780 428792 2786
rect 428740 2722 428792 2728
rect 427556 480 427584 2722
rect 428752 480 428780 2722
rect 429948 480 429976 5374
rect 430592 2854 430620 31010
rect 431880 26994 431908 40054
rect 431868 26988 431920 26994
rect 431868 26930 431920 26936
rect 432328 3460 432380 3466
rect 432328 3402 432380 3408
rect 430580 2848 430632 2854
rect 430580 2790 430632 2796
rect 431132 2780 431184 2786
rect 431132 2722 431184 2728
rect 431144 480 431172 2722
rect 432340 480 432368 3402
rect 433168 2922 433196 40054
rect 433260 39370 433288 43302
rect 433248 39364 433300 39370
rect 433248 39306 433300 39312
rect 433340 32496 433392 32502
rect 433340 32438 433392 32444
rect 433352 7682 433380 32438
rect 434640 28286 434668 43302
rect 434812 40928 434864 40934
rect 434812 40870 434864 40876
rect 434824 38622 434852 40870
rect 434812 38616 434864 38622
rect 434812 38558 434864 38564
rect 434812 29028 434864 29034
rect 434812 28970 434864 28976
rect 434628 28280 434680 28286
rect 434628 28222 434680 28228
rect 434824 19310 434852 28970
rect 434812 19304 434864 19310
rect 434812 19246 434864 19252
rect 434812 9784 434864 9790
rect 434812 9726 434864 9732
rect 434824 9654 434852 9726
rect 434812 9648 434864 9654
rect 434812 9590 434864 9596
rect 433340 7676 433392 7682
rect 433340 7618 433392 7624
rect 434628 7676 434680 7682
rect 434628 7618 434680 7624
rect 433522 4856 433578 4865
rect 433522 4791 433578 4800
rect 433156 2916 433208 2922
rect 433156 2858 433208 2864
rect 433536 480 433564 4791
rect 434640 480 434668 7618
rect 436020 3466 436048 43302
rect 437400 10334 437428 43302
rect 437952 40118 437980 43316
rect 439148 40118 439176 43316
rect 440344 40118 440372 43316
rect 441448 43302 441554 43330
rect 442750 43302 442948 43330
rect 443946 43302 444328 43330
rect 445142 43302 445708 43330
rect 437940 40112 437992 40118
rect 437940 40054 437992 40060
rect 438768 40112 438820 40118
rect 438768 40054 438820 40060
rect 439136 40112 439188 40118
rect 439136 40054 439188 40060
rect 440148 40112 440200 40118
rect 440148 40054 440200 40060
rect 440332 40112 440384 40118
rect 440332 40054 440384 40060
rect 438780 29646 438808 40054
rect 438768 29640 438820 29646
rect 438768 29582 438820 29588
rect 437480 28348 437532 28354
rect 437480 28290 437532 28296
rect 437388 10328 437440 10334
rect 437388 10270 437440 10276
rect 437020 5228 437072 5234
rect 437020 5170 437072 5176
rect 436008 3460 436060 3466
rect 436008 3402 436060 3408
rect 435824 604 435876 610
rect 435824 546 435876 552
rect 435836 480 435864 546
rect 437032 480 437060 5170
rect 437492 3346 437520 28290
rect 439412 4140 439464 4146
rect 439412 4082 439464 4088
rect 437492 3318 438256 3346
rect 438228 480 438256 3318
rect 439424 480 439452 4082
rect 440160 2990 440188 40054
rect 441448 31074 441476 43302
rect 441528 40112 441580 40118
rect 441528 40054 441580 40060
rect 441436 31068 441488 31074
rect 441436 31010 441488 31016
rect 441540 11830 441568 40054
rect 441528 11824 441580 11830
rect 441528 11766 441580 11772
rect 441620 11756 441672 11762
rect 441620 11698 441672 11704
rect 440608 5500 440660 5506
rect 440608 5442 440660 5448
rect 440148 2984 440200 2990
rect 440148 2926 440200 2932
rect 440620 480 440648 5442
rect 441632 3346 441660 11698
rect 442920 4146 442948 43302
rect 443184 40860 443236 40866
rect 443184 40802 443236 40808
rect 442908 4140 442960 4146
rect 442908 4082 442960 4088
rect 443196 3346 443224 40802
rect 444300 13190 444328 43302
rect 444380 33856 444432 33862
rect 444380 33798 444432 33804
rect 444288 13184 444340 13190
rect 444288 13126 444340 13132
rect 444196 4956 444248 4962
rect 444196 4898 444248 4904
rect 441632 3318 441844 3346
rect 441816 480 441844 3318
rect 443012 3318 443224 3346
rect 443012 480 443040 3318
rect 444208 480 444236 4898
rect 444392 3346 444420 33798
rect 445680 32502 445708 43302
rect 446232 40118 446260 43316
rect 447428 40118 447456 43316
rect 448624 40118 448652 43316
rect 446220 40112 446272 40118
rect 446220 40054 446272 40060
rect 447048 40112 447100 40118
rect 447048 40054 447100 40060
rect 447416 40112 447468 40118
rect 447416 40054 447468 40060
rect 448428 40112 448480 40118
rect 448428 40054 448480 40060
rect 448612 40112 448664 40118
rect 448612 40054 448664 40060
rect 449716 40112 449768 40118
rect 449716 40054 449768 40060
rect 445668 32496 445720 32502
rect 445668 32438 445720 32444
rect 446588 4004 446640 4010
rect 446588 3946 446640 3952
rect 444392 3318 445432 3346
rect 445404 480 445432 3318
rect 446600 480 446628 3946
rect 447060 3806 447088 40054
rect 448440 14482 448468 40054
rect 449728 33862 449756 40054
rect 449716 33856 449768 33862
rect 449716 33798 449768 33804
rect 448428 14476 448480 14482
rect 448428 14418 448480 14424
rect 448520 13116 448572 13122
rect 448520 13058 448572 13064
rect 447784 5296 447836 5302
rect 447784 5238 447836 5244
rect 447048 3800 447100 3806
rect 447048 3742 447100 3748
rect 447796 480 447824 5238
rect 448532 3346 448560 13058
rect 449820 3505 449848 43316
rect 449992 40792 450044 40798
rect 449992 40734 450044 40740
rect 449806 3496 449862 3505
rect 449806 3431 449862 3440
rect 450004 3346 450032 40734
rect 451016 37942 451044 43316
rect 452226 43302 452608 43330
rect 453422 43302 453988 43330
rect 454618 43302 455368 43330
rect 451004 37936 451056 37942
rect 451004 37878 451056 37884
rect 451280 35284 451332 35290
rect 451280 35226 451332 35232
rect 451292 3398 451320 35226
rect 452580 17270 452608 43302
rect 452568 17264 452620 17270
rect 452568 17206 452620 17212
rect 451372 4752 451424 4758
rect 451372 4694 451424 4700
rect 451280 3392 451332 3398
rect 448532 3318 449020 3346
rect 450004 3318 450216 3346
rect 451280 3334 451332 3340
rect 448992 480 449020 3318
rect 450188 480 450216 3318
rect 451384 2666 451412 4694
rect 453672 3936 453724 3942
rect 453672 3878 453724 3884
rect 452476 3392 452528 3398
rect 452476 3334 452528 3340
rect 451292 2638 451412 2666
rect 451292 480 451320 2638
rect 452488 480 452516 3334
rect 453684 480 453712 3878
rect 453960 3194 453988 43302
rect 455340 5438 455368 43302
rect 455800 40118 455828 43316
rect 456892 41132 456944 41138
rect 456892 41074 456944 41080
rect 455788 40112 455840 40118
rect 455788 40054 455840 40060
rect 456708 40112 456760 40118
rect 456708 40054 456760 40060
rect 456720 20058 456748 40054
rect 456708 20052 456760 20058
rect 456708 19994 456760 20000
rect 455420 14544 455472 14550
rect 455420 14486 455472 14492
rect 455328 5432 455380 5438
rect 455328 5374 455380 5380
rect 454868 5092 454920 5098
rect 454868 5034 454920 5040
rect 453948 3188 454000 3194
rect 453948 3130 454000 3136
rect 454880 480 454908 5034
rect 455432 610 455460 14486
rect 456904 610 456932 41074
rect 456996 40118 457024 43316
rect 458192 40118 458220 43316
rect 459388 40798 459416 43316
rect 460598 43302 460888 43330
rect 461794 43302 462268 43330
rect 462990 43302 463648 43330
rect 459376 40792 459428 40798
rect 459376 40734 459428 40740
rect 456984 40112 457036 40118
rect 456984 40054 457036 40060
rect 458088 40112 458140 40118
rect 458088 40054 458140 40060
rect 458180 40112 458232 40118
rect 458180 40054 458232 40060
rect 459468 40112 459520 40118
rect 459468 40054 459520 40060
rect 458100 3126 458128 40054
rect 458180 15904 458232 15910
rect 458180 15846 458232 15852
rect 458088 3120 458140 3126
rect 458088 3062 458140 3068
rect 458192 626 458220 15846
rect 459480 5370 459508 40054
rect 459652 6180 459704 6186
rect 459652 6122 459704 6128
rect 459468 5364 459520 5370
rect 459468 5306 459520 5312
rect 455420 604 455472 610
rect 455420 546 455472 552
rect 456064 604 456116 610
rect 456064 546 456116 552
rect 456892 604 456944 610
rect 456892 546 456944 552
rect 457260 604 457312 610
rect 458192 598 458496 626
rect 457260 546 457312 552
rect 456076 480 456104 546
rect 457272 480 457300 546
rect 458468 480 458496 598
rect 459664 480 459692 6122
rect 460756 3868 460808 3874
rect 460756 3810 460808 3816
rect 460768 3074 460796 3810
rect 460860 3262 460888 43302
rect 460940 17332 460992 17338
rect 460940 17274 460992 17280
rect 460952 3346 460980 17274
rect 462240 5302 462268 43302
rect 462320 38072 462372 38078
rect 462320 38014 462372 38020
rect 462228 5296 462280 5302
rect 462228 5238 462280 5244
rect 462332 3346 462360 38014
rect 463620 4962 463648 43302
rect 463792 41064 463844 41070
rect 463792 41006 463844 41012
rect 463608 4956 463660 4962
rect 463608 4898 463660 4904
rect 463804 3346 463832 41006
rect 464172 40118 464200 43316
rect 465368 40118 465396 43316
rect 466564 40118 466592 43316
rect 467104 40792 467156 40798
rect 467104 40734 467156 40740
rect 464160 40112 464212 40118
rect 464160 40054 464212 40060
rect 464988 40112 465040 40118
rect 464988 40054 465040 40060
rect 465356 40112 465408 40118
rect 465356 40054 465408 40060
rect 466368 40112 466420 40118
rect 466368 40054 466420 40060
rect 466552 40112 466604 40118
rect 466552 40054 466604 40060
rect 460952 3318 462084 3346
rect 462332 3318 463280 3346
rect 463804 3318 464476 3346
rect 460848 3256 460900 3262
rect 460848 3198 460900 3204
rect 460768 3046 460888 3074
rect 460860 480 460888 3046
rect 462056 480 462084 3318
rect 463252 480 463280 3318
rect 464448 480 464476 3318
rect 465000 3058 465028 40054
rect 465080 19984 465132 19990
rect 465080 19926 465132 19932
rect 464988 3052 465040 3058
rect 464988 2994 465040 3000
rect 465092 1714 465120 19926
rect 466380 5234 466408 40054
rect 466460 29708 466512 29714
rect 466460 29650 466512 29656
rect 466368 5228 466420 5234
rect 466368 5170 466420 5176
rect 466472 3346 466500 29650
rect 467116 18698 467144 40734
rect 467760 40730 467788 43316
rect 468970 43302 469168 43330
rect 470166 43302 470548 43330
rect 471362 43302 471928 43330
rect 467748 40724 467800 40730
rect 467748 40666 467800 40672
rect 467748 40112 467800 40118
rect 467748 40054 467800 40060
rect 467760 22846 467788 40054
rect 467748 22840 467800 22846
rect 467748 22782 467800 22788
rect 467104 18692 467156 18698
rect 467104 18634 467156 18640
rect 467840 18624 467892 18630
rect 467840 18566 467892 18572
rect 467852 3398 467880 18566
rect 469140 15910 469168 43302
rect 469220 26920 469272 26926
rect 469220 26862 469272 26868
rect 469128 15904 469180 15910
rect 469128 15846 469180 15852
rect 467840 3392 467892 3398
rect 466472 3318 466868 3346
rect 469128 3392 469180 3398
rect 467840 3334 467892 3340
rect 467930 3360 467986 3369
rect 465092 1686 465672 1714
rect 465644 480 465672 1686
rect 466840 480 466868 3318
rect 469128 3334 469180 3340
rect 469232 3346 469260 26862
rect 470520 21418 470548 43302
rect 470508 21412 470560 21418
rect 470508 21354 470560 21360
rect 471520 4072 471572 4078
rect 471520 4014 471572 4020
rect 467930 3295 467986 3304
rect 467944 480 467972 3295
rect 469140 480 469168 3334
rect 469232 3318 470364 3346
rect 470336 480 470364 3318
rect 471532 480 471560 4014
rect 471900 3398 471928 43302
rect 472452 40118 472480 43316
rect 473648 40118 473676 43316
rect 474844 40934 474872 43316
rect 474832 40928 474884 40934
rect 474832 40870 474884 40876
rect 472440 40112 472492 40118
rect 472440 40054 472492 40060
rect 473268 40112 473320 40118
rect 473268 40054 473320 40060
rect 473636 40112 473688 40118
rect 473636 40054 473688 40060
rect 474648 40112 474700 40118
rect 474648 40054 474700 40060
rect 471980 22772 472032 22778
rect 471980 22714 472032 22720
rect 471888 3392 471940 3398
rect 471888 3334 471940 3340
rect 471992 610 472020 22714
rect 473280 5166 473308 40054
rect 473360 35216 473412 35222
rect 473360 35158 473412 35164
rect 473268 5160 473320 5166
rect 473268 5102 473320 5108
rect 473372 610 473400 35158
rect 474660 24206 474688 40054
rect 474648 24200 474700 24206
rect 474648 24142 474700 24148
rect 476040 4826 476068 43316
rect 477250 43302 477448 43330
rect 478446 43302 478828 43330
rect 479642 43302 480208 43330
rect 476120 36576 476172 36582
rect 476120 36518 476172 36524
rect 476028 4820 476080 4826
rect 476028 4762 476080 4768
rect 475108 3596 475160 3602
rect 475108 3538 475160 3544
rect 471980 604 472032 610
rect 471980 546 472032 552
rect 472716 604 472768 610
rect 472716 546 472768 552
rect 473360 604 473412 610
rect 473360 546 473412 552
rect 473912 604 473964 610
rect 473912 546 473964 552
rect 472728 480 472756 546
rect 473924 480 473952 546
rect 475120 480 475148 3538
rect 476132 626 476160 36518
rect 477420 25566 477448 43302
rect 477408 25560 477460 25566
rect 477408 25502 477460 25508
rect 477592 10396 477644 10402
rect 477592 10338 477644 10344
rect 477604 626 477632 10338
rect 478696 3664 478748 3670
rect 478696 3606 478748 3612
rect 476132 598 476344 626
rect 476316 480 476344 598
rect 477512 598 477632 626
rect 477512 480 477540 598
rect 478708 480 478736 3606
rect 478800 3330 478828 43302
rect 478880 21480 478932 21486
rect 478880 21422 478932 21428
rect 478788 3324 478840 3330
rect 478788 3266 478840 3272
rect 478892 610 478920 21422
rect 480180 5098 480208 43302
rect 480824 40118 480852 43316
rect 482020 40798 482048 43316
rect 482008 40792 482060 40798
rect 482008 40734 482060 40740
rect 483216 40118 483244 43316
rect 484412 40118 484440 43316
rect 485622 43302 485728 43330
rect 486818 43302 487108 43330
rect 488014 43302 488488 43330
rect 480812 40112 480864 40118
rect 480812 40054 480864 40060
rect 481548 40112 481600 40118
rect 481548 40054 481600 40060
rect 483204 40112 483256 40118
rect 483204 40054 483256 40060
rect 484308 40112 484360 40118
rect 484308 40054 484360 40060
rect 484400 40112 484452 40118
rect 484400 40054 484452 40060
rect 485596 40112 485648 40118
rect 485596 40054 485648 40060
rect 480260 32428 480312 32434
rect 480260 32370 480312 32376
rect 480168 5092 480220 5098
rect 480168 5034 480220 5040
rect 480272 3482 480300 32370
rect 481560 7682 481588 40054
rect 481548 7676 481600 7682
rect 481548 7618 481600 7624
rect 483480 6248 483532 6254
rect 483480 6190 483532 6196
rect 482284 3732 482336 3738
rect 482284 3674 482336 3680
rect 480272 3454 481128 3482
rect 478880 604 478932 610
rect 478880 546 478932 552
rect 479892 604 479944 610
rect 479892 546 479944 552
rect 479904 480 479932 546
rect 481100 480 481128 3454
rect 482296 480 482324 3674
rect 483492 480 483520 6190
rect 484320 5030 484348 40054
rect 485608 26926 485636 40054
rect 485596 26920 485648 26926
rect 485596 26862 485648 26868
rect 484400 24132 484452 24138
rect 484400 24074 484452 24080
rect 484308 5024 484360 5030
rect 484308 4966 484360 4972
rect 484412 3482 484440 24074
rect 485700 3641 485728 43302
rect 485780 15972 485832 15978
rect 485780 15914 485832 15920
rect 485686 3632 485742 3641
rect 485686 3567 485742 3576
rect 484412 3454 484624 3482
rect 484596 480 484624 3454
rect 485792 480 485820 15914
rect 486976 7608 487028 7614
rect 486976 7550 487028 7556
rect 486988 480 487016 7550
rect 487080 4894 487108 43302
rect 488460 28354 488488 43302
rect 489196 40866 489224 43316
rect 489184 40860 489236 40866
rect 489184 40802 489236 40808
rect 490392 40118 490420 43316
rect 491588 40118 491616 43316
rect 492784 40118 492812 43316
rect 493888 43302 493994 43330
rect 495190 43302 495388 43330
rect 496386 43302 496768 43330
rect 497490 43302 498148 43330
rect 490380 40112 490432 40118
rect 490380 40054 490432 40060
rect 491208 40112 491260 40118
rect 491208 40054 491260 40060
rect 491576 40112 491628 40118
rect 491576 40054 491628 40060
rect 492588 40112 492640 40118
rect 492588 40054 492640 40060
rect 492772 40112 492824 40118
rect 492772 40054 492824 40060
rect 488448 28348 488500 28354
rect 488448 28290 488500 28296
rect 487160 25628 487212 25634
rect 487160 25570 487212 25576
rect 487068 4888 487120 4894
rect 487068 4830 487120 4836
rect 487172 3482 487200 25570
rect 491220 8974 491248 40054
rect 492600 31142 492628 40054
rect 493888 36582 493916 43302
rect 493968 40112 494020 40118
rect 493968 40054 494020 40060
rect 493876 36576 493928 36582
rect 493876 36518 493928 36524
rect 492588 31136 492640 31142
rect 492588 31078 492640 31084
rect 491300 26988 491352 26994
rect 491300 26930 491352 26936
rect 490564 8968 490616 8974
rect 490564 8910 490616 8916
rect 491208 8968 491260 8974
rect 491208 8910 491260 8916
rect 489368 3528 489420 3534
rect 487172 3454 488212 3482
rect 489368 3470 489420 3476
rect 488184 480 488212 3454
rect 489380 480 489408 3470
rect 490576 480 490604 8910
rect 491312 3482 491340 26930
rect 493980 4078 494008 40054
rect 494060 39364 494112 39370
rect 494060 39306 494112 39312
rect 493968 4072 494020 4078
rect 493968 4014 494020 4020
rect 494072 3482 494100 39306
rect 495360 32434 495388 43302
rect 495348 32428 495400 32434
rect 495348 32370 495400 32376
rect 494152 28280 494204 28286
rect 494152 28222 494204 28228
rect 494164 3602 494192 28222
rect 496740 4010 496768 43302
rect 498120 10334 498148 43302
rect 498672 40118 498700 43316
rect 499868 40118 499896 43316
rect 498660 40112 498712 40118
rect 498660 40054 498712 40060
rect 499488 40112 499540 40118
rect 499488 40054 499540 40060
rect 499856 40112 499908 40118
rect 499856 40054 499908 40060
rect 500868 40112 500920 40118
rect 500868 40054 500920 40060
rect 498200 29640 498252 29646
rect 498200 29582 498252 29588
rect 496820 10328 496872 10334
rect 496820 10270 496872 10276
rect 498108 10328 498160 10334
rect 498108 10270 498160 10276
rect 496728 4004 496780 4010
rect 496728 3946 496780 3952
rect 494152 3596 494204 3602
rect 494152 3538 494204 3544
rect 495348 3596 495400 3602
rect 495348 3538 495400 3544
rect 491312 3454 491800 3482
rect 494072 3454 494192 3482
rect 491772 480 491800 3454
rect 492956 2916 493008 2922
rect 492956 2858 493008 2864
rect 492968 480 492996 2858
rect 494164 480 494192 3454
rect 495360 480 495388 3538
rect 496832 3482 496860 10270
rect 498212 3482 498240 29582
rect 499500 11762 499528 40054
rect 499488 11756 499540 11762
rect 499488 11698 499540 11704
rect 500880 3942 500908 40054
rect 501064 39370 501092 43316
rect 502168 43302 502274 43330
rect 503470 43302 503668 43330
rect 504666 43302 505048 43330
rect 505862 43302 506428 43330
rect 507058 43302 507808 43330
rect 501052 39364 501104 39370
rect 501052 39306 501104 39312
rect 502168 33794 502196 43302
rect 502156 33788 502208 33794
rect 502156 33730 502208 33736
rect 502432 31068 502484 31074
rect 502432 31010 502484 31016
rect 500960 11824 501012 11830
rect 500960 11766 501012 11772
rect 500868 3936 500920 3942
rect 500868 3878 500920 3884
rect 500972 3482 501000 11766
rect 496544 3460 496596 3466
rect 496832 3454 497780 3482
rect 498212 3454 498976 3482
rect 500972 3454 501276 3482
rect 496544 3402 496596 3408
rect 496556 480 496584 3402
rect 497752 480 497780 3454
rect 498948 480 498976 3454
rect 500132 2984 500184 2990
rect 500132 2926 500184 2932
rect 500144 480 500172 2926
rect 501248 480 501276 3454
rect 502444 480 502472 31010
rect 503640 6882 503668 43302
rect 503720 13184 503772 13190
rect 503720 13126 503772 13132
rect 503456 6854 503668 6882
rect 503456 3874 503484 6854
rect 503628 4140 503680 4146
rect 503628 4082 503680 4088
rect 503444 3868 503496 3874
rect 503444 3810 503496 3816
rect 503640 480 503668 4082
rect 503732 3482 503760 13126
rect 505020 13122 505048 43302
rect 505100 32496 505152 32502
rect 505100 32438 505152 32444
rect 505008 13116 505060 13122
rect 505008 13058 505060 13064
rect 505112 3482 505140 32438
rect 506400 19990 506428 43302
rect 506388 19984 506440 19990
rect 506388 19926 506440 19932
rect 507216 3800 507268 3806
rect 507216 3742 507268 3748
rect 503732 3454 504864 3482
rect 505112 3454 506060 3482
rect 504836 480 504864 3454
rect 506032 480 506060 3454
rect 507228 480 507256 3742
rect 507780 3670 507808 43302
rect 508240 40118 508268 43316
rect 509436 40118 509464 43316
rect 510632 40118 510660 43316
rect 508228 40112 508280 40118
rect 508228 40054 508280 40060
rect 509148 40112 509200 40118
rect 509148 40054 509200 40060
rect 509424 40112 509476 40118
rect 509424 40054 509476 40060
rect 510528 40112 510580 40118
rect 510528 40054 510580 40060
rect 510620 40112 510672 40118
rect 510620 40054 510672 40060
rect 509160 14482 509188 40054
rect 509240 33856 509292 33862
rect 509240 33798 509292 33804
rect 507860 14476 507912 14482
rect 507860 14418 507912 14424
rect 509148 14476 509200 14482
rect 509148 14418 509200 14424
rect 507768 3664 507820 3670
rect 507768 3606 507820 3612
rect 507872 3482 507900 14418
rect 507872 3454 508452 3482
rect 508424 480 508452 3454
rect 509252 3346 509280 33798
rect 510540 18630 510568 40054
rect 511828 35222 511856 43316
rect 513038 43302 513328 43330
rect 514234 43302 514708 43330
rect 515430 43302 516088 43330
rect 511908 40112 511960 40118
rect 511908 40054 511960 40060
rect 511816 35216 511868 35222
rect 511816 35158 511868 35164
rect 510528 18624 510580 18630
rect 510528 18566 510580 18572
rect 511920 3738 511948 40054
rect 512000 37936 512052 37942
rect 512000 37878 512052 37884
rect 511908 3732 511960 3738
rect 511908 3674 511960 3680
rect 510802 3496 510858 3505
rect 510802 3431 510858 3440
rect 509252 3318 509648 3346
rect 509620 480 509648 3318
rect 510816 480 510844 3431
rect 512012 480 512040 37878
rect 512092 17264 512144 17270
rect 512092 17206 512144 17212
rect 512104 3346 512132 17206
rect 513300 3806 513328 43302
rect 514680 4146 514708 43302
rect 516060 6186 516088 43302
rect 516612 40118 516640 43316
rect 517808 40118 517836 43316
rect 516600 40112 516652 40118
rect 516600 40054 516652 40060
rect 517428 40112 517480 40118
rect 517428 40054 517480 40060
rect 517796 40112 517848 40118
rect 517796 40054 517848 40060
rect 518808 40112 518860 40118
rect 518808 40054 518860 40060
rect 516140 20052 516192 20058
rect 516140 19994 516192 20000
rect 516048 6180 516100 6186
rect 516048 6122 516100 6128
rect 515588 5432 515640 5438
rect 515588 5374 515640 5380
rect 514668 4140 514720 4146
rect 514668 4082 514720 4088
rect 513288 3800 513340 3806
rect 513288 3742 513340 3748
rect 512104 3318 513236 3346
rect 513208 480 513236 3318
rect 514392 3188 514444 3194
rect 514392 3130 514444 3136
rect 514404 480 514432 3130
rect 515600 480 515628 5374
rect 516152 3346 516180 19994
rect 517440 3602 517468 40054
rect 517428 3596 517480 3602
rect 517428 3538 517480 3544
rect 518820 3534 518848 40054
rect 519004 37942 519032 43316
rect 518992 37936 519044 37942
rect 518992 37878 519044 37884
rect 519084 5364 519136 5370
rect 519084 5306 519136 5312
rect 518808 3528 518860 3534
rect 518808 3470 518860 3476
rect 516152 3318 516824 3346
rect 516796 480 516824 3318
rect 517888 3120 517940 3126
rect 517888 3062 517940 3068
rect 517900 480 517928 3062
rect 519096 480 519124 5306
rect 520200 3369 520228 43316
rect 521410 43302 521608 43330
rect 520372 18692 520424 18698
rect 520372 18634 520424 18640
rect 520384 3482 520412 18634
rect 520292 3454 520412 3482
rect 521580 3466 521608 43302
rect 523696 41410 523724 76599
rect 523880 64870 523908 89927
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 523868 64864 523920 64870
rect 523868 64806 523920 64812
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 523866 63336 523922 63345
rect 523866 63271 523922 63280
rect 523774 50008 523830 50017
rect 523774 49943 523830 49952
rect 523684 41404 523736 41410
rect 523684 41346 523736 41352
rect 523788 17950 523816 49943
rect 523880 30326 523908 63271
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 535460 40928 535512 40934
rect 535460 40870 535512 40876
rect 528560 40724 528612 40730
rect 528560 40666 528612 40672
rect 523868 30320 523920 30326
rect 523868 30262 523920 30268
rect 527180 22840 527232 22846
rect 527180 22782 527232 22788
rect 523776 17944 523828 17950
rect 523776 17886 523828 17892
rect 522672 5296 522724 5302
rect 522672 5238 522724 5244
rect 521568 3460 521620 3466
rect 520186 3360 520242 3369
rect 520186 3295 520242 3304
rect 520292 480 520320 3454
rect 521568 3402 521620 3408
rect 521476 3256 521528 3262
rect 521476 3198 521528 3204
rect 521488 480 521516 3198
rect 522684 480 522712 5238
rect 526260 5228 526312 5234
rect 526260 5170 526312 5176
rect 523868 4956 523920 4962
rect 523868 4898 523920 4904
rect 523880 480 523908 4898
rect 525064 3052 525116 3058
rect 525064 2994 525116 3000
rect 525076 480 525104 2994
rect 526272 480 526300 5170
rect 527192 3346 527220 22782
rect 528572 3482 528600 40666
rect 534080 24200 534132 24206
rect 534080 24142 534132 24148
rect 529940 21412 529992 21418
rect 529940 21354 529992 21360
rect 528652 15904 528704 15910
rect 528652 15846 528704 15852
rect 528664 4214 528692 15846
rect 528652 4208 528704 4214
rect 528652 4150 528704 4156
rect 529848 4208 529900 4214
rect 529848 4150 529900 4156
rect 528572 3454 528692 3482
rect 527192 3318 527496 3346
rect 527468 480 527496 3318
rect 528664 480 528692 3454
rect 529860 480 529888 4150
rect 529952 3482 529980 21354
rect 533436 5160 533488 5166
rect 533436 5102 533488 5108
rect 529952 3454 531084 3482
rect 531056 480 531084 3454
rect 532240 3392 532292 3398
rect 532240 3334 532292 3340
rect 532252 480 532280 3334
rect 533448 480 533476 5102
rect 534092 3482 534120 24142
rect 535472 3482 535500 40870
rect 549260 40860 549312 40866
rect 549260 40802 549312 40808
rect 542360 40792 542412 40798
rect 542360 40734 542412 40740
rect 536840 25560 536892 25566
rect 536840 25502 536892 25508
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536852 3398 536880 25502
rect 541716 7676 541768 7682
rect 541716 7618 541768 7624
rect 540520 5092 540572 5098
rect 540520 5034 540572 5040
rect 536932 4820 536984 4826
rect 536932 4762 536984 4768
rect 536840 3392 536892 3398
rect 536840 3334 536892 3340
rect 536944 480 536972 4762
rect 538128 3392 538180 3398
rect 538128 3334 538180 3340
rect 538140 480 538168 3334
rect 539324 3324 539376 3330
rect 539324 3266 539376 3272
rect 539336 480 539364 3266
rect 540532 480 540560 5034
rect 541728 480 541756 7618
rect 542372 3482 542400 40734
rect 547880 28348 547932 28354
rect 547880 28290 547932 28296
rect 545120 26920 545172 26926
rect 545120 26862 545172 26868
rect 544108 5024 544160 5030
rect 544108 4966 544160 4972
rect 542372 3454 542952 3482
rect 542924 480 542952 3454
rect 544120 480 544148 4966
rect 545132 3482 545160 26862
rect 547696 4888 547748 4894
rect 547696 4830 547748 4836
rect 546498 3632 546554 3641
rect 546498 3567 546554 3576
rect 545132 3454 545344 3482
rect 545316 480 545344 3454
rect 546512 480 546540 3567
rect 547708 480 547736 4830
rect 547892 3482 547920 28290
rect 549272 3482 549300 40802
rect 561680 39364 561732 39370
rect 561680 39306 561732 39312
rect 554780 36576 554832 36582
rect 554780 36518 554832 36524
rect 552020 31136 552072 31142
rect 552020 31078 552072 31084
rect 551192 8968 551244 8974
rect 551192 8910 551244 8916
rect 547892 3454 548932 3482
rect 549272 3454 550128 3482
rect 548904 480 548932 3454
rect 550100 480 550128 3454
rect 551204 480 551232 8910
rect 552032 3482 552060 31078
rect 553584 4072 553636 4078
rect 553584 4014 553636 4020
rect 552032 3454 552428 3482
rect 552400 480 552428 3454
rect 553596 480 553624 4014
rect 554792 480 554820 36518
rect 554872 32428 554924 32434
rect 554872 32370 554924 32376
rect 554884 3482 554912 32370
rect 558920 11756 558972 11762
rect 558920 11698 558972 11704
rect 557540 10328 557592 10334
rect 557540 10270 557592 10276
rect 557172 4004 557224 4010
rect 557172 3946 557224 3952
rect 554884 3454 556016 3482
rect 555988 480 556016 3454
rect 557184 480 557212 3946
rect 557552 3482 557580 10270
rect 558932 3482 558960 11698
rect 560760 3936 560812 3942
rect 560760 3878 560812 3884
rect 557552 3454 558408 3482
rect 558932 3454 559604 3482
rect 558380 480 558408 3454
rect 559576 480 559604 3454
rect 560772 480 560800 3878
rect 561692 3482 561720 39306
rect 579620 37936 579672 37942
rect 579620 37878 579672 37884
rect 571432 35216 571484 35222
rect 571432 35158 571484 35164
rect 563152 33788 563204 33794
rect 563152 33730 563204 33736
rect 561692 3454 561996 3482
rect 561968 480 561996 3454
rect 563164 480 563192 33730
rect 565820 19984 565872 19990
rect 565820 19926 565872 19932
rect 564440 13116 564492 13122
rect 564440 13058 564492 13064
rect 564348 3868 564400 3874
rect 564348 3810 564400 3816
rect 564360 480 564388 3810
rect 564452 3482 564480 13058
rect 565832 3482 565860 19926
rect 569960 18624 570012 18630
rect 569960 18566 570012 18572
rect 568580 14476 568632 14482
rect 568580 14418 568632 14424
rect 567844 3664 567896 3670
rect 567844 3606 567896 3612
rect 564452 3454 565584 3482
rect 565832 3454 566780 3482
rect 565556 480 565584 3454
rect 566752 480 566780 3454
rect 567856 480 567884 3606
rect 568592 3482 568620 14418
rect 569972 3482 570000 18566
rect 571340 3732 571392 3738
rect 571340 3674 571392 3680
rect 568592 3454 569080 3482
rect 569972 3454 570276 3482
rect 569052 480 569080 3454
rect 570248 480 570276 3454
rect 571352 3210 571380 3674
rect 571444 3398 571472 35158
rect 576216 6180 576268 6186
rect 576216 6122 576268 6128
rect 575020 4140 575072 4146
rect 575020 4082 575072 4088
rect 573824 3800 573876 3806
rect 573824 3742 573876 3748
rect 571432 3392 571484 3398
rect 571432 3334 571484 3340
rect 572628 3392 572680 3398
rect 572628 3334 572680 3340
rect 571352 3182 571472 3210
rect 571444 480 571472 3182
rect 572640 480 572668 3334
rect 573836 480 573864 3742
rect 575032 480 575060 4082
rect 576228 480 576256 6122
rect 577412 3596 577464 3602
rect 577412 3538 577464 3544
rect 577424 480 577452 3538
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 578620 480 578648 3470
rect 579632 610 579660 37878
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 580080 17944 580132 17950
rect 580080 17886 580132 17892
rect 580092 17649 580120 17886
rect 580078 17640 580134 17649
rect 580078 17575 580134 17584
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 579620 604 579672 610
rect 579620 546 579672 552
rect 579804 604 579856 610
rect 579804 546 579856 552
rect 579816 480 579844 546
rect 581012 480 581040 3295
rect 582208 480 582236 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 682216 3478 682272
rect 3514 667936 3570 667992
rect 3422 624824 3478 624880
rect 3606 653520 3662 653576
rect 3514 610408 3570 610464
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 580170 697992 580226 698048
rect 59358 635976 59414 636032
rect 580170 686296 580226 686352
rect 580262 674600 580318 674656
rect 580170 639376 580226 639432
rect 523774 636520 523830 636576
rect 523682 623192 523738 623248
rect 59358 621696 59414 621752
rect 59358 607416 59414 607472
rect 523682 596536 523738 596592
rect 3606 595992 3662 596048
rect 3422 567296 3478 567352
rect 59358 593136 59414 593192
rect 59358 578856 59414 578912
rect 59358 564576 59414 564632
rect 3514 553016 3570 553072
rect 3422 538600 3478 538656
rect 59358 550296 59414 550352
rect 580446 651072 580502 651128
rect 580354 627680 580410 627736
rect 524326 609900 524328 609920
rect 524328 609900 524380 609920
rect 524380 609900 524382 609920
rect 524326 609864 524382 609900
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 523866 583208 523922 583264
rect 580262 580760 580318 580816
rect 524326 569900 524382 569936
rect 524326 569880 524328 569900
rect 524328 569880 524380 569900
rect 524380 569880 524382 569900
rect 580170 557232 580226 557288
rect 523774 556552 523830 556608
rect 523682 543224 523738 543280
rect 59358 536016 59414 536072
rect 523222 529896 523278 529952
rect 59358 521736 59414 521792
rect 3330 509904 3386 509960
rect 59358 507456 59414 507512
rect 580170 545536 580226 545592
rect 580354 533840 580410 533896
rect 523866 516568 523922 516624
rect 580170 510312 580226 510368
rect 523774 503240 523830 503296
rect 3330 495488 3386 495544
rect 59358 493176 59414 493232
rect 3606 481072 3662 481128
rect 59358 478896 59414 478952
rect 59358 464616 59414 464672
rect 3422 452376 3478 452432
rect 59358 450336 59414 450392
rect 580170 498616 580226 498672
rect 524326 489912 524382 489968
rect 580170 486784 580226 486840
rect 523866 476584 523922 476640
rect 580170 463392 580226 463448
rect 523774 463256 523830 463312
rect 523682 449928 523738 449984
rect 3422 437960 3478 438016
rect 59358 436092 59360 436112
rect 59360 436092 59412 436112
rect 59412 436092 59414 436112
rect 59358 436056 59414 436092
rect 3422 423680 3478 423736
rect 59358 421776 59414 421832
rect 580170 451696 580226 451752
rect 580170 439864 580226 439920
rect 523866 436600 523922 436656
rect 523774 423272 523830 423328
rect 580170 416472 580226 416528
rect 523682 409944 523738 410000
rect 59358 407496 59414 407552
rect 3514 394984 3570 395040
rect 59358 393216 59414 393272
rect 3422 380568 3478 380624
rect 59358 378936 59414 378992
rect 580170 404776 580226 404832
rect 523866 396616 523922 396672
rect 580170 392944 580226 393000
rect 523774 383288 523830 383344
rect 523682 369960 523738 370016
rect 580170 369552 580226 369608
rect 3514 366152 3570 366208
rect 59358 364656 59414 364712
rect 3422 337456 3478 337512
rect 580170 357856 580226 357912
rect 523682 356632 523738 356688
rect 59358 350376 59414 350432
rect 3514 323040 3570 323096
rect 3422 294344 3478 294400
rect 59358 335960 59414 336016
rect 580170 346024 580226 346080
rect 523774 343168 523830 343224
rect 523682 329840 523738 329896
rect 580170 322632 580226 322688
rect 59358 321680 59414 321736
rect 523498 316512 523554 316568
rect 579802 310800 579858 310856
rect 3606 308760 3662 308816
rect 59358 307400 59414 307456
rect 3514 280064 3570 280120
rect 523682 303184 523738 303240
rect 580170 299104 580226 299160
rect 59358 293120 59414 293176
rect 523222 289856 523278 289912
rect 59358 278840 59414 278896
rect 524326 276528 524382 276584
rect 580170 275712 580226 275768
rect 3698 265648 3754 265704
rect 59358 264560 59414 264616
rect 579802 263880 579858 263936
rect 3606 251232 3662 251288
rect 3422 236952 3478 237008
rect 3514 208120 3570 208176
rect 524326 263200 524382 263256
rect 580170 252184 580226 252240
rect 59358 250280 59414 250336
rect 523958 249872 524014 249928
rect 523682 236544 523738 236600
rect 59358 236020 59414 236056
rect 59358 236000 59360 236020
rect 59360 236000 59412 236020
rect 59412 236000 59414 236020
rect 580170 228792 580226 228848
rect 523682 223216 523738 223272
rect 3698 222536 3754 222592
rect 59358 221720 59414 221776
rect 580170 216960 580226 217016
rect 523406 209888 523462 209944
rect 59358 207440 59414 207496
rect 3606 193840 3662 193896
rect 3422 179424 3478 179480
rect 579802 205264 579858 205320
rect 523682 196560 523738 196616
rect 59358 193160 59414 193216
rect 523774 183232 523830 183288
rect 59358 178880 59414 178936
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 523682 169904 523738 169960
rect 3698 165008 3754 165064
rect 59358 164600 59414 164656
rect 579802 158344 579858 158400
rect 523682 156576 523738 156632
rect 3606 150728 3662 150784
rect 59358 150320 59414 150376
rect 3514 136312 3570 136368
rect 3422 122032 3478 122088
rect 59358 136040 59414 136096
rect 523866 143248 523922 143304
rect 523774 129920 523830 129976
rect 59358 121760 59414 121816
rect 523682 116592 523738 116648
rect 3698 107616 3754 107672
rect 59358 107480 59414 107536
rect 3606 93200 3662 93256
rect 3514 78920 3570 78976
rect 3422 35808 3478 35864
rect 59358 93200 59414 93256
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 523774 103264 523830 103320
rect 59358 78920 59414 78976
rect 523866 89936 523922 89992
rect 523682 76608 523738 76664
rect 59358 64640 59414 64696
rect 3790 64504 3846 64560
rect 59358 50360 59414 50416
rect 3698 50088 3754 50144
rect 3606 21392 3662 21448
rect 3514 7112 3570 7168
rect 85486 3440 85542 3496
rect 92294 3304 92350 3360
rect 146850 3440 146906 3496
rect 153934 3304 153990 3360
rect 339406 3304 339462 3360
rect 364246 3440 364302 3496
rect 383106 29008 383162 29064
rect 383290 29008 383346 29064
rect 390374 9696 390430 9752
rect 390650 9696 390706 9752
rect 400218 3304 400274 3360
rect 407026 3304 407082 3360
rect 425058 4820 425114 4856
rect 425058 4800 425060 4820
rect 425060 4800 425112 4820
rect 425112 4800 425114 4820
rect 425150 3440 425206 3496
rect 433522 4800 433578 4856
rect 449806 3440 449862 3496
rect 467930 3304 467986 3360
rect 485686 3576 485742 3632
rect 510802 3440 510858 3496
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 523866 63280 523922 63336
rect 523774 49952 523830 50008
rect 580170 40976 580226 41032
rect 520186 3304 520242 3360
rect 546498 3576 546554 3632
rect 580170 29280 580226 29336
rect 580078 17584 580134 17640
rect 580998 3304 581054 3360
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 3417 682274 3483 682277
rect -960 682272 3483 682274
rect -960 682216 3422 682272
rect 3478 682216 3483 682272
rect -960 682214 3483 682216
rect -960 682124 480 682214
rect 3417 682211 3483 682214
rect 580257 674658 580323 674661
rect 583520 674658 584960 674748
rect 580257 674656 584960 674658
rect 580257 674600 580262 674656
rect 580318 674600 584960 674656
rect 580257 674598 584960 674600
rect 580257 674595 580323 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3509 667994 3575 667997
rect -960 667992 3575 667994
rect -960 667936 3514 667992
rect 3570 667936 3575 667992
rect -960 667934 3575 667936
rect -960 667844 480 667934
rect 3509 667931 3575 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3601 653578 3667 653581
rect -960 653576 3667 653578
rect -960 653520 3606 653576
rect 3662 653520 3667 653576
rect -960 653518 3667 653520
rect -960 653428 480 653518
rect 3601 653515 3667 653518
rect 580441 651130 580507 651133
rect 583520 651130 584960 651220
rect 580441 651128 584960 651130
rect 580441 651072 580446 651128
rect 580502 651072 584960 651128
rect 580441 651070 584960 651072
rect 580441 651067 580507 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 523769 636578 523835 636581
rect 521916 636576 523835 636578
rect 521916 636520 523774 636576
rect 523830 636520 523835 636576
rect 521916 636518 523835 636520
rect 523769 636515 523835 636518
rect 59353 636034 59419 636037
rect 59353 636032 62100 636034
rect 59353 635976 59358 636032
rect 59414 635976 62100 636032
rect 59353 635974 62100 635976
rect 59353 635971 59419 635974
rect 580349 627738 580415 627741
rect 583520 627738 584960 627828
rect 580349 627736 584960 627738
rect 580349 627680 580354 627736
rect 580410 627680 584960 627736
rect 580349 627678 584960 627680
rect 580349 627675 580415 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 523677 623250 523743 623253
rect 521916 623248 523743 623250
rect 521916 623192 523682 623248
rect 523738 623192 523743 623248
rect 521916 623190 523743 623192
rect 523677 623187 523743 623190
rect 59353 621754 59419 621757
rect 59353 621752 62100 621754
rect 59353 621696 59358 621752
rect 59414 621696 62100 621752
rect 59353 621694 62100 621696
rect 59353 621691 59419 621694
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3509 610466 3575 610469
rect -960 610464 3575 610466
rect -960 610408 3514 610464
rect 3570 610408 3575 610464
rect -960 610406 3575 610408
rect -960 610316 480 610406
rect 3509 610403 3575 610406
rect 524321 609922 524387 609925
rect 521916 609920 524387 609922
rect 521916 609864 524326 609920
rect 524382 609864 524387 609920
rect 521916 609862 524387 609864
rect 524321 609859 524387 609862
rect 59353 607474 59419 607477
rect 59353 607472 62100 607474
rect 59353 607416 59358 607472
rect 59414 607416 62100 607472
rect 59353 607414 62100 607416
rect 59353 607411 59419 607414
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect 523677 596594 523743 596597
rect 521916 596592 523743 596594
rect 521916 596536 523682 596592
rect 523738 596536 523743 596592
rect 521916 596534 523743 596536
rect 523677 596531 523743 596534
rect -960 596050 480 596140
rect 3601 596050 3667 596053
rect -960 596048 3667 596050
rect -960 595992 3606 596048
rect 3662 595992 3667 596048
rect -960 595990 3667 595992
rect -960 595900 480 595990
rect 3601 595987 3667 595990
rect 59353 593194 59419 593197
rect 59353 593192 62100 593194
rect 59353 593136 59358 593192
rect 59414 593136 62100 593192
rect 59353 593134 62100 593136
rect 59353 593131 59419 593134
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect 523861 583266 523927 583269
rect 521916 583264 523927 583266
rect 521916 583208 523866 583264
rect 523922 583208 523927 583264
rect 521916 583206 523927 583208
rect 523861 583203 523927 583206
rect -960 581620 480 581860
rect 580257 580818 580323 580821
rect 583520 580818 584960 580908
rect 580257 580816 584960 580818
rect 580257 580760 580262 580816
rect 580318 580760 584960 580816
rect 580257 580758 584960 580760
rect 580257 580755 580323 580758
rect 583520 580668 584960 580758
rect 59353 578914 59419 578917
rect 59353 578912 62100 578914
rect 59353 578856 59358 578912
rect 59414 578856 62100 578912
rect 59353 578854 62100 578856
rect 59353 578851 59419 578854
rect 524321 569938 524387 569941
rect 521916 569936 524387 569938
rect 521916 569880 524326 569936
rect 524382 569880 524387 569936
rect 521916 569878 524387 569880
rect 524321 569875 524387 569878
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 59353 564634 59419 564637
rect 59353 564632 62100 564634
rect 59353 564576 59358 564632
rect 59414 564576 62100 564632
rect 59353 564574 62100 564576
rect 59353 564571 59419 564574
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect 523769 556610 523835 556613
rect 521916 556608 523835 556610
rect 521916 556552 523774 556608
rect 523830 556552 523835 556608
rect 521916 556550 523835 556552
rect 523769 556547 523835 556550
rect -960 553074 480 553164
rect 3509 553074 3575 553077
rect -960 553072 3575 553074
rect -960 553016 3514 553072
rect 3570 553016 3575 553072
rect -960 553014 3575 553016
rect -960 552924 480 553014
rect 3509 553011 3575 553014
rect 59353 550354 59419 550357
rect 59353 550352 62100 550354
rect 59353 550296 59358 550352
rect 59414 550296 62100 550352
rect 59353 550294 62100 550296
rect 59353 550291 59419 550294
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 523677 543282 523743 543285
rect 521916 543280 523743 543282
rect 521916 543224 523682 543280
rect 523738 543224 523743 543280
rect 521916 543222 523743 543224
rect 523677 543219 523743 543222
rect -960 538658 480 538748
rect 3417 538658 3483 538661
rect -960 538656 3483 538658
rect -960 538600 3422 538656
rect 3478 538600 3483 538656
rect -960 538598 3483 538600
rect -960 538508 480 538598
rect 3417 538595 3483 538598
rect 59353 536074 59419 536077
rect 59353 536072 62100 536074
rect 59353 536016 59358 536072
rect 59414 536016 62100 536072
rect 59353 536014 62100 536016
rect 59353 536011 59419 536014
rect 580349 533898 580415 533901
rect 583520 533898 584960 533988
rect 580349 533896 584960 533898
rect 580349 533840 580354 533896
rect 580410 533840 584960 533896
rect 580349 533838 584960 533840
rect 580349 533835 580415 533838
rect 583520 533748 584960 533838
rect 523217 529954 523283 529957
rect 521916 529952 523283 529954
rect 521916 529896 523222 529952
rect 523278 529896 523283 529952
rect 521916 529894 523283 529896
rect 523217 529891 523283 529894
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 59353 521794 59419 521797
rect 59353 521792 62100 521794
rect 59353 521736 59358 521792
rect 59414 521736 62100 521792
rect 59353 521734 62100 521736
rect 59353 521731 59419 521734
rect 523861 516626 523927 516629
rect 521916 516624 523927 516626
rect 521916 516568 523866 516624
rect 523922 516568 523927 516624
rect 521916 516566 523927 516568
rect 523861 516563 523927 516566
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3325 509962 3391 509965
rect -960 509960 3391 509962
rect -960 509904 3330 509960
rect 3386 509904 3391 509960
rect -960 509902 3391 509904
rect -960 509812 480 509902
rect 3325 509899 3391 509902
rect 59353 507514 59419 507517
rect 59353 507512 62100 507514
rect 59353 507456 59358 507512
rect 59414 507456 62100 507512
rect 59353 507454 62100 507456
rect 59353 507451 59419 507454
rect 523769 503298 523835 503301
rect 521916 503296 523835 503298
rect 521916 503240 523774 503296
rect 523830 503240 523835 503296
rect 521916 503238 523835 503240
rect 523769 503235 523835 503238
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 59353 493234 59419 493237
rect 59353 493232 62100 493234
rect 59353 493176 59358 493232
rect 59414 493176 62100 493232
rect 59353 493174 62100 493176
rect 59353 493171 59419 493174
rect 524321 489970 524387 489973
rect 521916 489968 524387 489970
rect 521916 489912 524326 489968
rect 524382 489912 524387 489968
rect 521916 489910 524387 489912
rect 524321 489907 524387 489910
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect -960 481130 480 481220
rect 3601 481130 3667 481133
rect -960 481128 3667 481130
rect -960 481072 3606 481128
rect 3662 481072 3667 481128
rect -960 481070 3667 481072
rect -960 480980 480 481070
rect 3601 481067 3667 481070
rect 59353 478954 59419 478957
rect 59353 478952 62100 478954
rect 59353 478896 59358 478952
rect 59414 478896 62100 478952
rect 59353 478894 62100 478896
rect 59353 478891 59419 478894
rect 523861 476642 523927 476645
rect 521916 476640 523927 476642
rect 521916 476584 523866 476640
rect 523922 476584 523927 476640
rect 521916 476582 523927 476584
rect 523861 476579 523927 476582
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 59353 464674 59419 464677
rect 59353 464672 62100 464674
rect 59353 464616 59358 464672
rect 59414 464616 62100 464672
rect 59353 464614 62100 464616
rect 59353 464611 59419 464614
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 523769 463314 523835 463317
rect 521916 463312 523835 463314
rect 521916 463256 523774 463312
rect 523830 463256 523835 463312
rect 583520 463300 584960 463390
rect 521916 463254 523835 463256
rect 523769 463251 523835 463254
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 59353 450394 59419 450397
rect 59353 450392 62100 450394
rect 59353 450336 59358 450392
rect 59414 450336 62100 450392
rect 59353 450334 62100 450336
rect 59353 450331 59419 450334
rect 523677 449986 523743 449989
rect 521916 449984 523743 449986
rect 521916 449928 523682 449984
rect 523738 449928 523743 449984
rect 521916 449926 523743 449928
rect 523677 449923 523743 449926
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3417 438018 3483 438021
rect -960 438016 3483 438018
rect -960 437960 3422 438016
rect 3478 437960 3483 438016
rect -960 437958 3483 437960
rect -960 437868 480 437958
rect 3417 437955 3483 437958
rect 523861 436658 523927 436661
rect 521916 436656 523927 436658
rect 521916 436600 523866 436656
rect 523922 436600 523927 436656
rect 521916 436598 523927 436600
rect 523861 436595 523927 436598
rect 59353 436114 59419 436117
rect 59353 436112 62100 436114
rect 59353 436056 59358 436112
rect 59414 436056 62100 436112
rect 59353 436054 62100 436056
rect 59353 436051 59419 436054
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3417 423738 3483 423741
rect -960 423736 3483 423738
rect -960 423680 3422 423736
rect 3478 423680 3483 423736
rect -960 423678 3483 423680
rect -960 423588 480 423678
rect 3417 423675 3483 423678
rect 523769 423330 523835 423333
rect 521916 423328 523835 423330
rect 521916 423272 523774 423328
rect 523830 423272 523835 423328
rect 521916 423270 523835 423272
rect 523769 423267 523835 423270
rect 59353 421834 59419 421837
rect 59353 421832 62100 421834
rect 59353 421776 59358 421832
rect 59414 421776 62100 421832
rect 59353 421774 62100 421776
rect 59353 421771 59419 421774
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect 523677 410002 523743 410005
rect 521916 410000 523743 410002
rect 521916 409944 523682 410000
rect 523738 409944 523743 410000
rect 521916 409942 523743 409944
rect 523677 409939 523743 409942
rect -960 409172 480 409412
rect 59353 407554 59419 407557
rect 59353 407552 62100 407554
rect 59353 407496 59358 407552
rect 59414 407496 62100 407552
rect 59353 407494 62100 407496
rect 59353 407491 59419 407494
rect 580165 404834 580231 404837
rect 583520 404834 584960 404924
rect 580165 404832 584960 404834
rect 580165 404776 580170 404832
rect 580226 404776 584960 404832
rect 580165 404774 584960 404776
rect 580165 404771 580231 404774
rect 583520 404684 584960 404774
rect 523861 396674 523927 396677
rect 521916 396672 523927 396674
rect 521916 396616 523866 396672
rect 523922 396616 523927 396672
rect 521916 396614 523927 396616
rect 523861 396611 523927 396614
rect -960 395042 480 395132
rect 3509 395042 3575 395045
rect -960 395040 3575 395042
rect -960 394984 3514 395040
rect 3570 394984 3575 395040
rect -960 394982 3575 394984
rect -960 394892 480 394982
rect 3509 394979 3575 394982
rect 59353 393274 59419 393277
rect 59353 393272 62100 393274
rect 59353 393216 59358 393272
rect 59414 393216 62100 393272
rect 59353 393214 62100 393216
rect 59353 393211 59419 393214
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 523769 383346 523835 383349
rect 521916 383344 523835 383346
rect 521916 383288 523774 383344
rect 523830 383288 523835 383344
rect 521916 383286 523835 383288
rect 523769 383283 523835 383286
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3417 380626 3483 380629
rect -960 380624 3483 380626
rect -960 380568 3422 380624
rect 3478 380568 3483 380624
rect -960 380566 3483 380568
rect -960 380476 480 380566
rect 3417 380563 3483 380566
rect 59353 378994 59419 378997
rect 59353 378992 62100 378994
rect 59353 378936 59358 378992
rect 59414 378936 62100 378992
rect 59353 378934 62100 378936
rect 59353 378931 59419 378934
rect 523677 370018 523743 370021
rect 521916 370016 523743 370018
rect 521916 369960 523682 370016
rect 523738 369960 523743 370016
rect 521916 369958 523743 369960
rect 523677 369955 523743 369958
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3509 366210 3575 366213
rect -960 366208 3575 366210
rect -960 366152 3514 366208
rect 3570 366152 3575 366208
rect -960 366150 3575 366152
rect -960 366060 480 366150
rect 3509 366147 3575 366150
rect 59353 364714 59419 364717
rect 59353 364712 62100 364714
rect 59353 364656 59358 364712
rect 59414 364656 62100 364712
rect 59353 364654 62100 364656
rect 59353 364651 59419 364654
rect 580165 357914 580231 357917
rect 583520 357914 584960 358004
rect 580165 357912 584960 357914
rect 580165 357856 580170 357912
rect 580226 357856 584960 357912
rect 580165 357854 584960 357856
rect 580165 357851 580231 357854
rect 583520 357764 584960 357854
rect 523677 356690 523743 356693
rect 521916 356688 523743 356690
rect 521916 356632 523682 356688
rect 523738 356632 523743 356688
rect 521916 356630 523743 356632
rect 523677 356627 523743 356630
rect -960 351780 480 352020
rect 59353 350434 59419 350437
rect 59353 350432 62100 350434
rect 59353 350376 59358 350432
rect 59414 350376 62100 350432
rect 59353 350374 62100 350376
rect 59353 350371 59419 350374
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 523769 343226 523835 343229
rect 521916 343224 523835 343226
rect 521916 343168 523774 343224
rect 523830 343168 523835 343224
rect 521916 343166 523835 343168
rect 523769 343163 523835 343166
rect -960 337514 480 337604
rect 3417 337514 3483 337517
rect -960 337512 3483 337514
rect -960 337456 3422 337512
rect 3478 337456 3483 337512
rect -960 337454 3483 337456
rect -960 337364 480 337454
rect 3417 337451 3483 337454
rect 59353 336018 59419 336021
rect 59353 336016 62100 336018
rect 59353 335960 59358 336016
rect 59414 335960 62100 336016
rect 59353 335958 62100 335960
rect 59353 335955 59419 335958
rect 583520 334236 584960 334476
rect 523677 329898 523743 329901
rect 521916 329896 523743 329898
rect 521916 329840 523682 329896
rect 523738 329840 523743 329896
rect 521916 329838 523743 329840
rect 523677 329835 523743 329838
rect -960 323098 480 323188
rect 3509 323098 3575 323101
rect -960 323096 3575 323098
rect -960 323040 3514 323096
rect 3570 323040 3575 323096
rect -960 323038 3575 323040
rect -960 322948 480 323038
rect 3509 323035 3575 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 59353 321738 59419 321741
rect 59353 321736 62100 321738
rect 59353 321680 59358 321736
rect 59414 321680 62100 321736
rect 59353 321678 62100 321680
rect 59353 321675 59419 321678
rect 523493 316570 523559 316573
rect 521916 316568 523559 316570
rect 521916 316512 523498 316568
rect 523554 316512 523559 316568
rect 521916 316510 523559 316512
rect 523493 316507 523559 316510
rect 579797 310858 579863 310861
rect 583520 310858 584960 310948
rect 579797 310856 584960 310858
rect 579797 310800 579802 310856
rect 579858 310800 584960 310856
rect 579797 310798 584960 310800
rect 579797 310795 579863 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3601 308818 3667 308821
rect -960 308816 3667 308818
rect -960 308760 3606 308816
rect 3662 308760 3667 308816
rect -960 308758 3667 308760
rect -960 308668 480 308758
rect 3601 308755 3667 308758
rect 59353 307458 59419 307461
rect 59353 307456 62100 307458
rect 59353 307400 59358 307456
rect 59414 307400 62100 307456
rect 59353 307398 62100 307400
rect 59353 307395 59419 307398
rect 523677 303242 523743 303245
rect 521916 303240 523743 303242
rect 521916 303184 523682 303240
rect 523738 303184 523743 303240
rect 521916 303182 523743 303184
rect 523677 303179 523743 303182
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3417 294402 3483 294405
rect -960 294400 3483 294402
rect -960 294344 3422 294400
rect 3478 294344 3483 294400
rect -960 294342 3483 294344
rect -960 294252 480 294342
rect 3417 294339 3483 294342
rect 59353 293178 59419 293181
rect 59353 293176 62100 293178
rect 59353 293120 59358 293176
rect 59414 293120 62100 293176
rect 59353 293118 62100 293120
rect 59353 293115 59419 293118
rect 523217 289914 523283 289917
rect 521916 289912 523283 289914
rect 521916 289856 523222 289912
rect 523278 289856 523283 289912
rect 521916 289854 523283 289856
rect 523217 289851 523283 289854
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3509 280122 3575 280125
rect -960 280120 3575 280122
rect -960 280064 3514 280120
rect 3570 280064 3575 280120
rect -960 280062 3575 280064
rect -960 279972 480 280062
rect 3509 280059 3575 280062
rect 59353 278898 59419 278901
rect 59353 278896 62100 278898
rect 59353 278840 59358 278896
rect 59414 278840 62100 278896
rect 59353 278838 62100 278840
rect 59353 278835 59419 278838
rect 524321 276586 524387 276589
rect 521916 276584 524387 276586
rect 521916 276528 524326 276584
rect 524382 276528 524387 276584
rect 521916 276526 524387 276528
rect 524321 276523 524387 276526
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect -960 265706 480 265796
rect 3693 265706 3759 265709
rect -960 265704 3759 265706
rect -960 265648 3698 265704
rect 3754 265648 3759 265704
rect -960 265646 3759 265648
rect -960 265556 480 265646
rect 3693 265643 3759 265646
rect 59353 264618 59419 264621
rect 59353 264616 62100 264618
rect 59353 264560 59358 264616
rect 59414 264560 62100 264616
rect 59353 264558 62100 264560
rect 59353 264555 59419 264558
rect 579797 263938 579863 263941
rect 583520 263938 584960 264028
rect 579797 263936 584960 263938
rect 579797 263880 579802 263936
rect 579858 263880 584960 263936
rect 579797 263878 584960 263880
rect 579797 263875 579863 263878
rect 583520 263788 584960 263878
rect 524321 263258 524387 263261
rect 521916 263256 524387 263258
rect 521916 263200 524326 263256
rect 524382 263200 524387 263256
rect 521916 263198 524387 263200
rect 524321 263195 524387 263198
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3601 251290 3667 251293
rect -960 251288 3667 251290
rect -960 251232 3606 251288
rect 3662 251232 3667 251288
rect -960 251230 3667 251232
rect -960 251140 480 251230
rect 3601 251227 3667 251230
rect 59353 250338 59419 250341
rect 59353 250336 62100 250338
rect 59353 250280 59358 250336
rect 59414 250280 62100 250336
rect 59353 250278 62100 250280
rect 59353 250275 59419 250278
rect 523953 249930 524019 249933
rect 521916 249928 524019 249930
rect 521916 249872 523958 249928
rect 524014 249872 524019 249928
rect 521916 249870 524019 249872
rect 523953 249867 524019 249870
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3417 237010 3483 237013
rect -960 237008 3483 237010
rect -960 236952 3422 237008
rect 3478 236952 3483 237008
rect -960 236950 3483 236952
rect -960 236860 480 236950
rect 3417 236947 3483 236950
rect 523677 236602 523743 236605
rect 521916 236600 523743 236602
rect 521916 236544 523682 236600
rect 523738 236544 523743 236600
rect 521916 236542 523743 236544
rect 523677 236539 523743 236542
rect 59353 236058 59419 236061
rect 59353 236056 62100 236058
rect 59353 236000 59358 236056
rect 59414 236000 62100 236056
rect 59353 235998 62100 236000
rect 59353 235995 59419 235998
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect 523677 223274 523743 223277
rect 521916 223272 523743 223274
rect 521916 223216 523682 223272
rect 523738 223216 523743 223272
rect 521916 223214 523743 223216
rect 523677 223211 523743 223214
rect -960 222594 480 222684
rect 3693 222594 3759 222597
rect -960 222592 3759 222594
rect -960 222536 3698 222592
rect 3754 222536 3759 222592
rect -960 222534 3759 222536
rect -960 222444 480 222534
rect 3693 222531 3759 222534
rect 59353 221778 59419 221781
rect 59353 221776 62100 221778
rect 59353 221720 59358 221776
rect 59414 221720 62100 221776
rect 59353 221718 62100 221720
rect 59353 221715 59419 221718
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 523401 209946 523467 209949
rect 521916 209944 523467 209946
rect 521916 209888 523406 209944
rect 523462 209888 523467 209944
rect 521916 209886 523467 209888
rect 523401 209883 523467 209886
rect -960 208178 480 208268
rect 3509 208178 3575 208181
rect -960 208176 3575 208178
rect -960 208120 3514 208176
rect 3570 208120 3575 208176
rect -960 208118 3575 208120
rect -960 208028 480 208118
rect 3509 208115 3575 208118
rect 59353 207498 59419 207501
rect 59353 207496 62100 207498
rect 59353 207440 59358 207496
rect 59414 207440 62100 207496
rect 59353 207438 62100 207440
rect 59353 207435 59419 207438
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 523677 196618 523743 196621
rect 521916 196616 523743 196618
rect 521916 196560 523682 196616
rect 523738 196560 523743 196616
rect 521916 196558 523743 196560
rect 523677 196555 523743 196558
rect -960 193898 480 193988
rect 3601 193898 3667 193901
rect -960 193896 3667 193898
rect -960 193840 3606 193896
rect 3662 193840 3667 193896
rect -960 193838 3667 193840
rect -960 193748 480 193838
rect 3601 193835 3667 193838
rect 583520 193476 584960 193716
rect 59353 193218 59419 193221
rect 59353 193216 62100 193218
rect 59353 193160 59358 193216
rect 59414 193160 62100 193216
rect 59353 193158 62100 193160
rect 59353 193155 59419 193158
rect 523769 183290 523835 183293
rect 521916 183288 523835 183290
rect 521916 183232 523774 183288
rect 523830 183232 523835 183288
rect 521916 183230 523835 183232
rect 523769 183227 523835 183230
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3417 179482 3483 179485
rect -960 179480 3483 179482
rect -960 179424 3422 179480
rect 3478 179424 3483 179480
rect -960 179422 3483 179424
rect -960 179332 480 179422
rect 3417 179419 3483 179422
rect 59353 178938 59419 178941
rect 59353 178936 62100 178938
rect 59353 178880 59358 178936
rect 59414 178880 62100 178936
rect 59353 178878 62100 178880
rect 59353 178875 59419 178878
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 523677 169962 523743 169965
rect 521916 169960 523743 169962
rect 521916 169904 523682 169960
rect 523738 169904 523743 169960
rect 583520 169948 584960 170038
rect 521916 169902 523743 169904
rect 523677 169899 523743 169902
rect -960 165066 480 165156
rect 3693 165066 3759 165069
rect -960 165064 3759 165066
rect -960 165008 3698 165064
rect 3754 165008 3759 165064
rect -960 165006 3759 165008
rect -960 164916 480 165006
rect 3693 165003 3759 165006
rect 59353 164658 59419 164661
rect 59353 164656 62100 164658
rect 59353 164600 59358 164656
rect 59414 164600 62100 164656
rect 59353 164598 62100 164600
rect 59353 164595 59419 164598
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 523677 156634 523743 156637
rect 521916 156632 523743 156634
rect 521916 156576 523682 156632
rect 523738 156576 523743 156632
rect 521916 156574 523743 156576
rect 523677 156571 523743 156574
rect -960 150786 480 150876
rect 3601 150786 3667 150789
rect -960 150784 3667 150786
rect -960 150728 3606 150784
rect 3662 150728 3667 150784
rect -960 150726 3667 150728
rect -960 150636 480 150726
rect 3601 150723 3667 150726
rect 59353 150378 59419 150381
rect 59353 150376 62100 150378
rect 59353 150320 59358 150376
rect 59414 150320 62100 150376
rect 59353 150318 62100 150320
rect 59353 150315 59419 150318
rect 583520 146556 584960 146796
rect 523861 143306 523927 143309
rect 521916 143304 523927 143306
rect 521916 143248 523866 143304
rect 523922 143248 523927 143304
rect 521916 143246 523927 143248
rect 523861 143243 523927 143246
rect -960 136370 480 136460
rect 3509 136370 3575 136373
rect -960 136368 3575 136370
rect -960 136312 3514 136368
rect 3570 136312 3575 136368
rect -960 136310 3575 136312
rect -960 136220 480 136310
rect 3509 136307 3575 136310
rect 59353 136098 59419 136101
rect 59353 136096 62100 136098
rect 59353 136040 59358 136096
rect 59414 136040 62100 136096
rect 59353 136038 62100 136040
rect 59353 136035 59419 136038
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 523769 129978 523835 129981
rect 521916 129976 523835 129978
rect 521916 129920 523774 129976
rect 523830 129920 523835 129976
rect 521916 129918 523835 129920
rect 523769 129915 523835 129918
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3417 122090 3483 122093
rect -960 122088 3483 122090
rect -960 122032 3422 122088
rect 3478 122032 3483 122088
rect -960 122030 3483 122032
rect -960 121940 480 122030
rect 3417 122027 3483 122030
rect 59353 121818 59419 121821
rect 59353 121816 62100 121818
rect 59353 121760 59358 121816
rect 59414 121760 62100 121816
rect 59353 121758 62100 121760
rect 59353 121755 59419 121758
rect 523677 116650 523743 116653
rect 521916 116648 523743 116650
rect 521916 116592 523682 116648
rect 523738 116592 523743 116648
rect 521916 116590 523743 116592
rect 523677 116587 523743 116590
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3693 107674 3759 107677
rect -960 107672 3759 107674
rect -960 107616 3698 107672
rect 3754 107616 3759 107672
rect -960 107614 3759 107616
rect -960 107524 480 107614
rect 3693 107611 3759 107614
rect 59353 107538 59419 107541
rect 59353 107536 62100 107538
rect 59353 107480 59358 107536
rect 59414 107480 62100 107536
rect 59353 107478 62100 107480
rect 59353 107475 59419 107478
rect 523769 103322 523835 103325
rect 521916 103320 523835 103322
rect 521916 103264 523774 103320
rect 523830 103264 523835 103320
rect 521916 103262 523835 103264
rect 523769 103259 523835 103262
rect 583520 99636 584960 99876
rect -960 93258 480 93348
rect 3601 93258 3667 93261
rect -960 93256 3667 93258
rect -960 93200 3606 93256
rect 3662 93200 3667 93256
rect -960 93198 3667 93200
rect -960 93108 480 93198
rect 3601 93195 3667 93198
rect 59353 93258 59419 93261
rect 59353 93256 62100 93258
rect 59353 93200 59358 93256
rect 59414 93200 62100 93256
rect 59353 93198 62100 93200
rect 59353 93195 59419 93198
rect 523861 89994 523927 89997
rect 521916 89992 523927 89994
rect 521916 89936 523866 89992
rect 523922 89936 523927 89992
rect 521916 89934 523927 89936
rect 523861 89931 523927 89934
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 3509 78978 3575 78981
rect -960 78976 3575 78978
rect -960 78920 3514 78976
rect 3570 78920 3575 78976
rect -960 78918 3575 78920
rect -960 78828 480 78918
rect 3509 78915 3575 78918
rect 59353 78978 59419 78981
rect 59353 78976 62100 78978
rect 59353 78920 59358 78976
rect 59414 78920 62100 78976
rect 59353 78918 62100 78920
rect 59353 78915 59419 78918
rect 523677 76666 523743 76669
rect 521916 76664 523743 76666
rect 521916 76608 523682 76664
rect 523738 76608 523743 76664
rect 521916 76606 523743 76608
rect 523677 76603 523743 76606
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 59353 64698 59419 64701
rect 59353 64696 62100 64698
rect -960 64562 480 64652
rect 59353 64640 59358 64696
rect 59414 64640 62100 64696
rect 59353 64638 62100 64640
rect 59353 64635 59419 64638
rect 3785 64562 3851 64565
rect -960 64560 3851 64562
rect -960 64504 3790 64560
rect 3846 64504 3851 64560
rect -960 64502 3851 64504
rect -960 64412 480 64502
rect 3785 64499 3851 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 523861 63338 523927 63341
rect 521916 63336 523927 63338
rect 521916 63280 523866 63336
rect 523922 63280 523927 63336
rect 521916 63278 523927 63280
rect 523861 63275 523927 63278
rect 583520 52716 584960 52956
rect 59353 50418 59419 50421
rect 59353 50416 62100 50418
rect 59353 50360 59358 50416
rect 59414 50360 62100 50416
rect 59353 50358 62100 50360
rect 59353 50355 59419 50358
rect -960 50146 480 50236
rect 3693 50146 3759 50149
rect -960 50144 3759 50146
rect -960 50088 3698 50144
rect 3754 50088 3759 50144
rect -960 50086 3759 50088
rect -960 49996 480 50086
rect 3693 50083 3759 50086
rect 523769 50010 523835 50013
rect 521916 50008 523835 50010
rect 521916 49952 523774 50008
rect 523830 49952 523835 50008
rect 521916 49950 523835 49952
rect 523769 49947 523835 49950
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect 383101 29066 383167 29069
rect 383285 29066 383351 29069
rect 383101 29064 383351 29066
rect 383101 29008 383106 29064
rect 383162 29008 383290 29064
rect 383346 29008 383351 29064
rect 383101 29006 383351 29008
rect 383101 29003 383167 29006
rect 383285 29003 383351 29006
rect -960 21450 480 21540
rect 3601 21450 3667 21453
rect -960 21448 3667 21450
rect -960 21392 3606 21448
rect 3662 21392 3667 21448
rect -960 21390 3667 21392
rect -960 21300 480 21390
rect 3601 21387 3667 21390
rect 580073 17642 580139 17645
rect 583520 17642 584960 17732
rect 580073 17640 584960 17642
rect 580073 17584 580078 17640
rect 580134 17584 584960 17640
rect 580073 17582 584960 17584
rect 580073 17579 580139 17582
rect 583520 17492 584960 17582
rect 390369 9754 390435 9757
rect 390645 9754 390711 9757
rect 390369 9752 390711 9754
rect 390369 9696 390374 9752
rect 390430 9696 390650 9752
rect 390706 9696 390711 9752
rect 390369 9694 390711 9696
rect 390369 9691 390435 9694
rect 390645 9691 390711 9694
rect -960 7170 480 7260
rect 3509 7170 3575 7173
rect -960 7168 3575 7170
rect -960 7112 3514 7168
rect 3570 7112 3575 7168
rect -960 7110 3575 7112
rect -960 7020 480 7110
rect 3509 7107 3575 7110
rect 583520 5796 584960 6036
rect 425053 4858 425119 4861
rect 433517 4858 433583 4861
rect 425053 4856 433583 4858
rect 425053 4800 425058 4856
rect 425114 4800 433522 4856
rect 433578 4800 433583 4856
rect 425053 4798 433583 4800
rect 425053 4795 425119 4798
rect 433517 4795 433583 4798
rect 485681 3634 485747 3637
rect 546493 3634 546559 3637
rect 485681 3632 546559 3634
rect 485681 3576 485686 3632
rect 485742 3576 546498 3632
rect 546554 3576 546559 3632
rect 485681 3574 546559 3576
rect 485681 3571 485747 3574
rect 546493 3571 546559 3574
rect 85481 3498 85547 3501
rect 146845 3498 146911 3501
rect 85481 3496 146911 3498
rect 85481 3440 85486 3496
rect 85542 3440 146850 3496
rect 146906 3440 146911 3496
rect 85481 3438 146911 3440
rect 85481 3435 85547 3438
rect 146845 3435 146911 3438
rect 364241 3498 364307 3501
rect 425145 3498 425211 3501
rect 364241 3496 425211 3498
rect 364241 3440 364246 3496
rect 364302 3440 425150 3496
rect 425206 3440 425211 3496
rect 364241 3438 425211 3440
rect 364241 3435 364307 3438
rect 425145 3435 425211 3438
rect 449801 3498 449867 3501
rect 510797 3498 510863 3501
rect 449801 3496 510863 3498
rect 449801 3440 449806 3496
rect 449862 3440 510802 3496
rect 510858 3440 510863 3496
rect 449801 3438 510863 3440
rect 449801 3435 449867 3438
rect 510797 3435 510863 3438
rect 92289 3362 92355 3365
rect 153929 3362 153995 3365
rect 92289 3360 153995 3362
rect 92289 3304 92294 3360
rect 92350 3304 153934 3360
rect 153990 3304 153995 3360
rect 92289 3302 153995 3304
rect 92289 3299 92355 3302
rect 153929 3299 153995 3302
rect 339401 3362 339467 3365
rect 400213 3362 400279 3365
rect 339401 3360 400279 3362
rect 339401 3304 339406 3360
rect 339462 3304 400218 3360
rect 400274 3304 400279 3360
rect 339401 3302 400279 3304
rect 339401 3299 339467 3302
rect 400213 3299 400279 3302
rect 407021 3362 407087 3365
rect 467925 3362 467991 3365
rect 407021 3360 467991 3362
rect 407021 3304 407026 3360
rect 407082 3304 467930 3360
rect 467986 3304 467991 3360
rect 407021 3302 467991 3304
rect 407021 3299 407087 3302
rect 467925 3299 467991 3302
rect 520181 3362 520247 3365
rect 580993 3362 581059 3365
rect 520181 3360 581059 3362
rect 520181 3304 520186 3360
rect 520242 3304 580998 3360
rect 581054 3304 581059 3360
rect 520181 3302 581059 3304
rect 520181 3299 520247 3302
rect 580993 3299 581059 3302
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 -6926 -7976 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 -5986 -7036 709922
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 -5046 -6096 708982
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 -4106 -5156 708042
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 -3166 -4216 707102
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 -2226 -3276 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 645200 73404 649898
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 645200 91404 667898
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 645200 109404 649898
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 645200 127404 667898
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 645200 145404 649898
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 645200 163404 667898
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 645200 181404 649898
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 645200 199404 667898
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 645200 217404 649898
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 645200 235404 667898
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 645200 253404 649898
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 645200 271404 667898
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 645200 289404 649898
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 645200 307404 667898
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 645200 325404 649898
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 645200 343404 667898
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 645200 361404 649898
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 645200 379404 667898
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 645200 397404 649898
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 645200 415404 667898
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 645200 433404 649898
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 645200 451404 667898
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 645200 469404 649898
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 645200 487404 667898
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 645200 505404 649898
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 645200 523404 667898
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 81568 632454 81888 632476
rect 81568 632218 81610 632454
rect 81846 632218 81888 632454
rect 81568 632134 81888 632218
rect 81568 631898 81610 632134
rect 81846 631898 81888 632134
rect 81568 631876 81888 631898
rect 66208 614454 66528 614476
rect 66208 614218 66250 614454
rect 66486 614218 66528 614454
rect 66208 614134 66528 614218
rect 66208 613898 66250 614134
rect 66486 613898 66528 614134
rect 66208 613876 66528 613898
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 81568 596454 81888 596476
rect 81568 596218 81610 596454
rect 81846 596218 81888 596454
rect 81568 596134 81888 596218
rect 81568 595898 81610 596134
rect 81846 595898 81888 596134
rect 81568 595876 81888 595898
rect 66208 578454 66528 578476
rect 66208 578218 66250 578454
rect 66486 578218 66528 578454
rect 66208 578134 66528 578218
rect 66208 577898 66250 578134
rect 66486 577898 66528 578134
rect 66208 577876 66528 577898
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 81568 560454 81888 560476
rect 81568 560218 81610 560454
rect 81846 560218 81888 560454
rect 81568 560134 81888 560218
rect 81568 559898 81610 560134
rect 81846 559898 81888 560134
rect 81568 559876 81888 559898
rect 66208 542454 66528 542476
rect 66208 542218 66250 542454
rect 66486 542218 66528 542454
rect 66208 542134 66528 542218
rect 66208 541898 66250 542134
rect 66486 541898 66528 542134
rect 66208 541876 66528 541898
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 81568 524454 81888 524476
rect 81568 524218 81610 524454
rect 81846 524218 81888 524454
rect 81568 524134 81888 524218
rect 81568 523898 81610 524134
rect 81846 523898 81888 524134
rect 81568 523876 81888 523898
rect 66208 506454 66528 506476
rect 66208 506218 66250 506454
rect 66486 506218 66528 506454
rect 66208 506134 66528 506218
rect 66208 505898 66250 506134
rect 66486 505898 66528 506134
rect 66208 505876 66528 505898
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 81568 488454 81888 488476
rect 81568 488218 81610 488454
rect 81846 488218 81888 488454
rect 81568 488134 81888 488218
rect 81568 487898 81610 488134
rect 81846 487898 81888 488134
rect 81568 487876 81888 487898
rect 66208 470454 66528 470476
rect 66208 470218 66250 470454
rect 66486 470218 66528 470454
rect 66208 470134 66528 470218
rect 66208 469898 66250 470134
rect 66486 469898 66528 470134
rect 66208 469876 66528 469898
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 81568 452454 81888 452476
rect 81568 452218 81610 452454
rect 81846 452218 81888 452454
rect 81568 452134 81888 452218
rect 81568 451898 81610 452134
rect 81846 451898 81888 452134
rect 81568 451876 81888 451898
rect 66208 434454 66528 434476
rect 66208 434218 66250 434454
rect 66486 434218 66528 434454
rect 66208 434134 66528 434218
rect 66208 433898 66250 434134
rect 66486 433898 66528 434134
rect 66208 433876 66528 433898
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 81568 416454 81888 416476
rect 81568 416218 81610 416454
rect 81846 416218 81888 416454
rect 81568 416134 81888 416218
rect 81568 415898 81610 416134
rect 81846 415898 81888 416134
rect 81568 415876 81888 415898
rect 66208 398454 66528 398476
rect 66208 398218 66250 398454
rect 66486 398218 66528 398454
rect 66208 398134 66528 398218
rect 66208 397898 66250 398134
rect 66486 397898 66528 398134
rect 66208 397876 66528 397898
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 81568 380454 81888 380476
rect 81568 380218 81610 380454
rect 81846 380218 81888 380454
rect 81568 380134 81888 380218
rect 81568 379898 81610 380134
rect 81846 379898 81888 380134
rect 81568 379876 81888 379898
rect 66208 362454 66528 362476
rect 66208 362218 66250 362454
rect 66486 362218 66528 362454
rect 66208 362134 66528 362218
rect 66208 361898 66250 362134
rect 66486 361898 66528 362134
rect 66208 361876 66528 361898
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 81568 344454 81888 344476
rect 81568 344218 81610 344454
rect 81846 344218 81888 344454
rect 81568 344134 81888 344218
rect 81568 343898 81610 344134
rect 81846 343898 81888 344134
rect 81568 343876 81888 343898
rect 66208 326454 66528 326476
rect 66208 326218 66250 326454
rect 66486 326218 66528 326454
rect 66208 326134 66528 326218
rect 66208 325898 66250 326134
rect 66486 325898 66528 326134
rect 66208 325876 66528 325898
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 81568 308454 81888 308476
rect 81568 308218 81610 308454
rect 81846 308218 81888 308454
rect 81568 308134 81888 308218
rect 81568 307898 81610 308134
rect 81846 307898 81888 308134
rect 81568 307876 81888 307898
rect 66208 290454 66528 290476
rect 66208 290218 66250 290454
rect 66486 290218 66528 290454
rect 66208 290134 66528 290218
rect 66208 289898 66250 290134
rect 66486 289898 66528 290134
rect 66208 289876 66528 289898
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 81568 272454 81888 272476
rect 81568 272218 81610 272454
rect 81846 272218 81888 272454
rect 81568 272134 81888 272218
rect 81568 271898 81610 272134
rect 81846 271898 81888 272134
rect 81568 271876 81888 271898
rect 66208 254454 66528 254476
rect 66208 254218 66250 254454
rect 66486 254218 66528 254454
rect 66208 254134 66528 254218
rect 66208 253898 66250 254134
rect 66486 253898 66528 254134
rect 66208 253876 66528 253898
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 81568 236454 81888 236476
rect 81568 236218 81610 236454
rect 81846 236218 81888 236454
rect 81568 236134 81888 236218
rect 81568 235898 81610 236134
rect 81846 235898 81888 236134
rect 81568 235876 81888 235898
rect 66208 218454 66528 218476
rect 66208 218218 66250 218454
rect 66486 218218 66528 218454
rect 66208 218134 66528 218218
rect 66208 217898 66250 218134
rect 66486 217898 66528 218134
rect 66208 217876 66528 217898
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 81568 200454 81888 200476
rect 81568 200218 81610 200454
rect 81846 200218 81888 200454
rect 81568 200134 81888 200218
rect 81568 199898 81610 200134
rect 81846 199898 81888 200134
rect 81568 199876 81888 199898
rect 66208 182454 66528 182476
rect 66208 182218 66250 182454
rect 66486 182218 66528 182454
rect 66208 182134 66528 182218
rect 66208 181898 66250 182134
rect 66486 181898 66528 182134
rect 66208 181876 66528 181898
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 81568 164454 81888 164476
rect 81568 164218 81610 164454
rect 81846 164218 81888 164454
rect 81568 164134 81888 164218
rect 81568 163898 81610 164134
rect 81846 163898 81888 164134
rect 81568 163876 81888 163898
rect 66208 146454 66528 146476
rect 66208 146218 66250 146454
rect 66486 146218 66528 146454
rect 66208 146134 66528 146218
rect 66208 145898 66250 146134
rect 66486 145898 66528 146134
rect 66208 145876 66528 145898
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 81568 128454 81888 128476
rect 81568 128218 81610 128454
rect 81846 128218 81888 128454
rect 81568 128134 81888 128218
rect 81568 127898 81610 128134
rect 81846 127898 81888 128134
rect 81568 127876 81888 127898
rect 66208 110454 66528 110476
rect 66208 110218 66250 110454
rect 66486 110218 66528 110454
rect 66208 110134 66528 110218
rect 66208 109898 66250 110134
rect 66486 109898 66528 110134
rect 66208 109876 66528 109898
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 81568 92454 81888 92476
rect 81568 92218 81610 92454
rect 81846 92218 81888 92454
rect 81568 92134 81888 92218
rect 81568 91898 81610 92134
rect 81846 91898 81888 92134
rect 81568 91876 81888 91898
rect 66208 74454 66528 74476
rect 66208 74218 66250 74454
rect 66486 74218 66528 74454
rect 66208 74134 66528 74218
rect 66208 73898 66250 74134
rect 66486 73898 66528 74134
rect 66208 73876 66528 73898
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 81568 56454 81888 56476
rect 81568 56218 81610 56454
rect 81846 56218 81888 56454
rect 81568 56134 81888 56218
rect 81568 55898 81610 56134
rect 81846 55898 81888 56134
rect 81568 55876 81888 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 72804 38454 73404 41200
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 90804 20454 91404 41200
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 108804 38454 109404 41200
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 126804 20454 127404 41200
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 144804 38454 145404 41200
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 162804 20454 163404 41200
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 180804 38454 181404 41200
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 198804 20454 199404 41200
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 216804 38454 217404 41200
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 234804 20454 235404 41200
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 252804 38454 253404 41200
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 270804 20454 271404 41200
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 288804 38454 289404 41200
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 306804 20454 307404 41200
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 324804 38454 325404 41200
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 342804 20454 343404 41200
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 360804 38454 361404 41200
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 378804 20454 379404 41200
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 396804 38454 397404 41200
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 414804 20454 415404 41200
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 432804 38454 433404 41200
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 450804 20454 451404 41200
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 468804 38454 469404 41200
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 486804 20454 487404 41200
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 504804 38454 505404 41200
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 522804 20454 523404 41200
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 576804 704838 577404 705800
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 587200 -2226 587800 706162
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 588140 -3166 588740 707102
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 589080 -4106 589680 708042
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 590020 -5046 590620 708982
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 590960 -5986 591560 709922
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 591900 -6926 592500 710862
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 81610 632218 81846 632454
rect 81610 631898 81846 632134
rect 66250 614218 66486 614454
rect 66250 613898 66486 614134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 81610 596218 81846 596454
rect 81610 595898 81846 596134
rect 66250 578218 66486 578454
rect 66250 577898 66486 578134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 81610 560218 81846 560454
rect 81610 559898 81846 560134
rect 66250 542218 66486 542454
rect 66250 541898 66486 542134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 81610 524218 81846 524454
rect 81610 523898 81846 524134
rect 66250 506218 66486 506454
rect 66250 505898 66486 506134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 81610 488218 81846 488454
rect 81610 487898 81846 488134
rect 66250 470218 66486 470454
rect 66250 469898 66486 470134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 81610 452218 81846 452454
rect 81610 451898 81846 452134
rect 66250 434218 66486 434454
rect 66250 433898 66486 434134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 81610 416218 81846 416454
rect 81610 415898 81846 416134
rect 66250 398218 66486 398454
rect 66250 397898 66486 398134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 81610 380218 81846 380454
rect 81610 379898 81846 380134
rect 66250 362218 66486 362454
rect 66250 361898 66486 362134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 81610 344218 81846 344454
rect 81610 343898 81846 344134
rect 66250 326218 66486 326454
rect 66250 325898 66486 326134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 81610 308218 81846 308454
rect 81610 307898 81846 308134
rect 66250 290218 66486 290454
rect 66250 289898 66486 290134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 81610 272218 81846 272454
rect 81610 271898 81846 272134
rect 66250 254218 66486 254454
rect 66250 253898 66486 254134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 81610 236218 81846 236454
rect 81610 235898 81846 236134
rect 66250 218218 66486 218454
rect 66250 217898 66486 218134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 81610 200218 81846 200454
rect 81610 199898 81846 200134
rect 66250 182218 66486 182454
rect 66250 181898 66486 182134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 81610 164218 81846 164454
rect 81610 163898 81846 164134
rect 66250 146218 66486 146454
rect 66250 145898 66486 146134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 81610 128218 81846 128454
rect 81610 127898 81846 128134
rect 66250 110218 66486 110454
rect 66250 109898 66486 110134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 81610 92218 81846 92454
rect 81610 91898 81846 92134
rect 66250 74218 66486 74454
rect 66250 73898 66486 74134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 81610 56218 81846 56454
rect 81610 55898 81846 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 81568 632476 81888 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 81610 632454
rect 81846 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 81610 632134
rect 81846 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 81568 631874 81888 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 66208 614476 66528 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 66250 614454
rect 66486 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 66250 614134
rect 66486 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 66208 613874 66528 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 81568 596476 81888 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 81610 596454
rect 81846 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 81610 596134
rect 81846 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 81568 595874 81888 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 66208 578476 66528 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 66250 578454
rect 66486 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 66250 578134
rect 66486 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 66208 577874 66528 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 81568 560476 81888 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 81610 560454
rect 81846 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 81610 560134
rect 81846 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 81568 559874 81888 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 66208 542476 66528 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 66250 542454
rect 66486 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 66250 542134
rect 66486 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 66208 541874 66528 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 81568 524476 81888 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 81610 524454
rect 81846 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 81610 524134
rect 81846 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 81568 523874 81888 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 66208 506476 66528 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 66250 506454
rect 66486 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 66250 506134
rect 66486 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 66208 505874 66528 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 81568 488476 81888 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 81610 488454
rect 81846 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 81610 488134
rect 81846 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 81568 487874 81888 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 66208 470476 66528 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 66250 470454
rect 66486 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 66250 470134
rect 66486 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 66208 469874 66528 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 81568 452476 81888 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 81610 452454
rect 81846 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 81610 452134
rect 81846 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 81568 451874 81888 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 66208 434476 66528 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 66250 434454
rect 66486 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 66250 434134
rect 66486 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 66208 433874 66528 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 81568 416476 81888 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 81610 416454
rect 81846 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 81610 416134
rect 81846 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 81568 415874 81888 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 66208 398476 66528 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 66250 398454
rect 66486 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 66250 398134
rect 66486 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 66208 397874 66528 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 81568 380476 81888 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 81610 380454
rect 81846 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 81610 380134
rect 81846 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 81568 379874 81888 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 66208 362476 66528 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 66250 362454
rect 66486 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 66250 362134
rect 66486 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 66208 361874 66528 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 81568 344476 81888 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 81610 344454
rect 81846 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 81610 344134
rect 81846 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 81568 343874 81888 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 66208 326476 66528 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 66250 326454
rect 66486 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 66250 326134
rect 66486 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 66208 325874 66528 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 81568 308476 81888 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 81610 308454
rect 81846 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 81610 308134
rect 81846 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 81568 307874 81888 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 66208 290476 66528 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 66250 290454
rect 66486 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 66250 290134
rect 66486 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 66208 289874 66528 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 81568 272476 81888 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 81610 272454
rect 81846 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 81610 272134
rect 81846 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 81568 271874 81888 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 66208 254476 66528 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 66250 254454
rect 66486 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 66250 254134
rect 66486 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 66208 253874 66528 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 81568 236476 81888 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 81610 236454
rect 81846 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 81610 236134
rect 81846 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 81568 235874 81888 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 66208 218476 66528 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 66250 218454
rect 66486 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 66250 218134
rect 66486 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 66208 217874 66528 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 81568 200476 81888 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 81610 200454
rect 81846 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 81610 200134
rect 81846 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 81568 199874 81888 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 66208 182476 66528 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 66250 182454
rect 66486 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 66250 182134
rect 66486 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 66208 181874 66528 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 81568 164476 81888 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 81610 164454
rect 81846 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 81610 164134
rect 81846 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 81568 163874 81888 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 66208 146476 66528 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 66250 146454
rect 66486 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 66250 146134
rect 66486 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 66208 145874 66528 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 81568 128476 81888 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 81610 128454
rect 81846 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 81610 128134
rect 81846 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 81568 127874 81888 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 66208 110476 66528 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 66250 110454
rect 66486 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 66250 110134
rect 66486 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 66208 109874 66528 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 81568 92476 81888 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 81610 92454
rect 81846 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 81610 92134
rect 81846 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 81568 91874 81888 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 66208 74476 66528 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 66250 74454
rect 66486 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 66250 74134
rect 66486 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 66208 73874 66528 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 81568 56476 81888 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 81610 56454
rect 81846 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 81610 56134
rect 81846 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 81568 55874 81888 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 591900 -7506 592500 -7504
use ghazi_top_dffram_csv  mprj
timestamp 1609742308
transform 1 0 62000 0 1 43200
box 0 0 460000 600000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew signal input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew signal input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew signal input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew signal input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew signal input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew signal input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew signal input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew signal input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew signal input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew signal input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew signal input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew signal input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew signal input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew signal input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew signal input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew signal input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew signal input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew signal input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew signal input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew signal input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew signal input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew signal input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew signal input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew signal input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew signal input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew signal input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew signal input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew signal input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew signal input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew signal tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew signal tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew signal tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew signal tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew signal tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew signal tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew signal tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew signal tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew signal tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew signal tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew signal tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew signal tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew signal tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew signal tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew signal tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew signal tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew signal tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew signal tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew signal tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew signal tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew signal tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew signal tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew signal tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew signal tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew signal tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew signal tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew signal tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew signal tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew signal tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew signal tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew signal tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew signal tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew signal tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew signal tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew signal tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew signal tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew signal tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew signal tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew signal tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew signal tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew signal tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew signal tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew signal tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew signal tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew signal tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew signal tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew signal tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew signal tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew signal tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew signal tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew signal tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew signal tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew signal tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew signal tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew signal tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew signal tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew signal tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew signal tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew signal tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew signal tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew signal tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew signal tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew signal tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew signal tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew signal tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew signal tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew signal tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew signal tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew signal tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew signal tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew signal tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew signal tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew signal tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew signal tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew signal tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew signal tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew signal tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew signal tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew signal tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew signal tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew signal tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew signal tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew signal tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew signal tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew signal tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew signal tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew signal tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew signal tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew signal tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew signal tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew signal tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew signal tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew signal tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew signal tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew signal tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew signal tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew signal tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew signal tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew signal tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew signal tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew signal tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew signal tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew signal tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew signal tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew signal tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew signal tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew signal tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew signal tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew signal tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew signal tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew signal tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew signal tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew signal tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew signal tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew signal tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew signal tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew signal tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew signal tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew signal tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew signal tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew signal tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew signal tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew signal tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew signal tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew signal tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew signal tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew signal tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew signal tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew signal tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew signal tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew signal tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew signal tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew signal tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew signal tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew signal tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew signal tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew signal tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew signal tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew signal tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew signal tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew signal tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew signal tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew signal tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew signal tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew signal tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew signal tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew signal tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew signal tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew signal tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew signal tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew signal tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew signal tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew signal tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew signal tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew signal tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew signal tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew signal tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew signal tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew signal tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew signal tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew signal tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew signal tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew signal tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew signal tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew signal tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew signal tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew signal tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew signal tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew signal tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew signal tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew signal tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew signal tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew signal tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew signal tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew signal tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew signal tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew signal tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew signal tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew signal tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew signal tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew signal tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew signal tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew signal tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew signal tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew signal tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew signal input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew signal input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew signal input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew signal input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew signal input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew signal input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew signal input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew signal input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew signal input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew signal input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew signal input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew signal input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew signal input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew signal input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew signal input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew signal input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew signal input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew signal input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew signal input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew signal input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew signal input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew signal input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew signal input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew signal input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew signal input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew signal input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew signal input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew signal input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew signal input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew signal input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew signal input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew signal input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew signal input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew signal input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew signal input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew signal input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew signal input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew signal input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew signal input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew signal input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew signal input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew signal input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew signal input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew signal input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew signal input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew signal input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew signal input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew signal input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew signal input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew signal input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew signal input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew signal input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew signal input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew signal input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew signal input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew signal input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew signal input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew signal input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew signal input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew signal input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew signal input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew signal input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew signal input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew signal input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew signal input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew signal input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew signal input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew signal input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew signal input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew signal input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew signal input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew signal input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew signal input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew signal input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew signal input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew signal input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew signal input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew signal input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew signal input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew signal input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew signal input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew signal input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew signal input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew signal input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew signal input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew signal input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew signal input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew signal input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew signal input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew signal input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew signal input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew signal input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew signal input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew signal input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew signal input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew signal input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew signal input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew signal input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew signal input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew signal input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew signal input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew signal input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew signal input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew signal input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew signal input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew signal input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew signal input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew signal input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew signal input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew signal input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew signal input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew signal input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew signal input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew signal input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew signal input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew signal input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew signal input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew signal input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew signal input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew signal input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew signal input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew signal input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew signal input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew signal input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew signal input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew signal input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew signal input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew signal input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew signal input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew signal input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew signal input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew signal input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew signal input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew signal input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew signal input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew signal input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew signal input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew signal input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew signal input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew signal input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew signal input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew signal input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew signal input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew signal input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew signal input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew signal input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew signal input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew signal input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew signal input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew signal input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew signal input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew signal input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew signal input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew signal input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew signal input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew signal input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew signal input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew signal input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew signal input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew signal input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew signal input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew signal input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew signal input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew signal input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew signal input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew signal input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew signal input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew signal input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew signal input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew signal input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew signal input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew signal input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew signal input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew signal input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew signal input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew signal input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew signal input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew signal input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew signal input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew signal input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew signal input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew signal input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew signal input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew signal input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew signal input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew signal input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew signal input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew signal input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew signal tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew signal tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew signal tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew signal tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew signal tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew signal tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew signal tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew signal tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew signal tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew signal tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew signal tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew signal tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew signal tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew signal tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew signal tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew signal tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew signal tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew signal tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew signal tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew signal tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew signal tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew signal tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew signal tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew signal tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew signal tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew signal tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew signal tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew signal tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew signal tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew signal tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew signal tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew signal tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew signal input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew signal input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew signal input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew signal input
rlabel metal4 s 576804 -1864 577404 705800 6 vccd1
port 636 nsew power bidirectional
rlabel metal4 s 540804 -1864 541404 705800 6 vccd1.extra1
port 637 nsew power bidirectional
rlabel metal4 s 504804 645200 505404 705800 6 vccd1.extra2
port 638 nsew power bidirectional
rlabel metal4 s 468804 645200 469404 705800 6 vccd1.extra3
port 639 nsew power bidirectional
rlabel metal4 s 432804 645200 433404 705800 6 vccd1.extra4
port 640 nsew power bidirectional
rlabel metal4 s 396804 645200 397404 705800 6 vccd1.extra5
port 641 nsew power bidirectional
rlabel metal4 s 360804 645200 361404 705800 6 vccd1.extra6
port 642 nsew power bidirectional
rlabel metal4 s 324804 645200 325404 705800 6 vccd1.extra7
port 643 nsew power bidirectional
rlabel metal4 s 288804 645200 289404 705800 6 vccd1.extra8
port 644 nsew power bidirectional
rlabel metal4 s 252804 645200 253404 705800 6 vccd1.extra9
port 645 nsew power bidirectional
rlabel metal4 s 216804 645200 217404 705800 6 vccd1.extra10
port 646 nsew power bidirectional
rlabel metal4 s 180804 645200 181404 705800 6 vccd1.extra11
port 647 nsew power bidirectional
rlabel metal4 s 144804 645200 145404 705800 6 vccd1.extra12
port 648 nsew power bidirectional
rlabel metal4 s 108804 645200 109404 705800 6 vccd1.extra13
port 649 nsew power bidirectional
rlabel metal4 s 72804 645200 73404 705800 6 vccd1.extra14
port 650 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 705800 6 vccd1.extra15
port 651 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 705800 6 vccd1.extra16
port 652 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1.extra17
port 653 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1.extra18
port 654 nsew power bidirectional
rlabel metal4 s 504804 -1864 505404 41200 6 vccd1.extra19
port 655 nsew power bidirectional
rlabel metal4 s 468804 -1864 469404 41200 6 vccd1.extra20
port 656 nsew power bidirectional
rlabel metal4 s 432804 -1864 433404 41200 6 vccd1.extra21
port 657 nsew power bidirectional
rlabel metal4 s 396804 -1864 397404 41200 6 vccd1.extra22
port 658 nsew power bidirectional
rlabel metal4 s 360804 -1864 361404 41200 6 vccd1.extra23
port 659 nsew power bidirectional
rlabel metal4 s 324804 -1864 325404 41200 6 vccd1.extra24
port 660 nsew power bidirectional
rlabel metal4 s 288804 -1864 289404 41200 6 vccd1.extra25
port 661 nsew power bidirectional
rlabel metal4 s 252804 -1864 253404 41200 6 vccd1.extra26
port 662 nsew power bidirectional
rlabel metal4 s 216804 -1864 217404 41200 6 vccd1.extra27
port 663 nsew power bidirectional
rlabel metal4 s 180804 -1864 181404 41200 6 vccd1.extra28
port 664 nsew power bidirectional
rlabel metal4 s 144804 -1864 145404 41200 6 vccd1.extra29
port 665 nsew power bidirectional
rlabel metal4 s 108804 -1864 109404 41200 6 vccd1.extra30
port 666 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 41200 6 vccd1.extra31
port 667 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1.extra32
port 668 nsew power bidirectional
rlabel metal5 s -2936 685876 586860 686476 6 vccd1.extra33
port 669 nsew power bidirectional
rlabel metal5 s -2936 649876 586860 650476 6 vccd1.extra34
port 670 nsew power bidirectional
rlabel metal5 s -2936 613876 586860 614476 6 vccd1.extra35
port 671 nsew power bidirectional
rlabel metal5 s -2936 577876 586860 578476 6 vccd1.extra36
port 672 nsew power bidirectional
rlabel metal5 s -2936 541876 586860 542476 6 vccd1.extra37
port 673 nsew power bidirectional
rlabel metal5 s -2936 505876 586860 506476 6 vccd1.extra38
port 674 nsew power bidirectional
rlabel metal5 s -2936 469876 586860 470476 6 vccd1.extra39
port 675 nsew power bidirectional
rlabel metal5 s -2936 433876 586860 434476 6 vccd1.extra40
port 676 nsew power bidirectional
rlabel metal5 s -2936 397876 586860 398476 6 vccd1.extra41
port 677 nsew power bidirectional
rlabel metal5 s -2936 361876 586860 362476 6 vccd1.extra42
port 678 nsew power bidirectional
rlabel metal5 s -2936 325876 586860 326476 6 vccd1.extra43
port 679 nsew power bidirectional
rlabel metal5 s -2936 289876 586860 290476 6 vccd1.extra44
port 680 nsew power bidirectional
rlabel metal5 s -2936 253876 586860 254476 6 vccd1.extra45
port 681 nsew power bidirectional
rlabel metal5 s -2936 217876 586860 218476 6 vccd1.extra46
port 682 nsew power bidirectional
rlabel metal5 s -2936 181876 586860 182476 6 vccd1.extra47
port 683 nsew power bidirectional
rlabel metal5 s -2936 145876 586860 146476 6 vccd1.extra48
port 684 nsew power bidirectional
rlabel metal5 s -2936 109876 586860 110476 6 vccd1.extra49
port 685 nsew power bidirectional
rlabel metal5 s -2936 73876 586860 74476 6 vccd1.extra50
port 686 nsew power bidirectional
rlabel metal5 s -2936 37876 586860 38476 6 vccd1.extra51
port 687 nsew power bidirectional
rlabel metal5 s -2936 1876 586860 2476 6 vccd1.extra52
port 688 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1.extra53
port 689 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 690 nsew ground bidirectional
rlabel metal4 s 558804 -1864 559404 705800 6 vssd1.extra1
port 691 nsew ground bidirectional
rlabel metal4 s 522804 645200 523404 705800 6 vssd1.extra2
port 692 nsew ground bidirectional
rlabel metal4 s 486804 645200 487404 705800 6 vssd1.extra3
port 693 nsew ground bidirectional
rlabel metal4 s 450804 645200 451404 705800 6 vssd1.extra4
port 694 nsew ground bidirectional
rlabel metal4 s 414804 645200 415404 705800 6 vssd1.extra5
port 695 nsew ground bidirectional
rlabel metal4 s 378804 645200 379404 705800 6 vssd1.extra6
port 696 nsew ground bidirectional
rlabel metal4 s 342804 645200 343404 705800 6 vssd1.extra7
port 697 nsew ground bidirectional
rlabel metal4 s 306804 645200 307404 705800 6 vssd1.extra8
port 698 nsew ground bidirectional
rlabel metal4 s 270804 645200 271404 705800 6 vssd1.extra9
port 699 nsew ground bidirectional
rlabel metal4 s 234804 645200 235404 705800 6 vssd1.extra10
port 700 nsew ground bidirectional
rlabel metal4 s 198804 645200 199404 705800 6 vssd1.extra11
port 701 nsew ground bidirectional
rlabel metal4 s 162804 645200 163404 705800 6 vssd1.extra12
port 702 nsew ground bidirectional
rlabel metal4 s 126804 645200 127404 705800 6 vssd1.extra13
port 703 nsew ground bidirectional
rlabel metal4 s 90804 645200 91404 705800 6 vssd1.extra14
port 704 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 705800 6 vssd1.extra15
port 705 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 705800 6 vssd1.extra16
port 706 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1.extra17
port 707 nsew ground bidirectional
rlabel metal4 s 522804 -1864 523404 41200 6 vssd1.extra18
port 708 nsew ground bidirectional
rlabel metal4 s 486804 -1864 487404 41200 6 vssd1.extra19
port 709 nsew ground bidirectional
rlabel metal4 s 450804 -1864 451404 41200 6 vssd1.extra20
port 710 nsew ground bidirectional
rlabel metal4 s 414804 -1864 415404 41200 6 vssd1.extra21
port 711 nsew ground bidirectional
rlabel metal4 s 378804 -1864 379404 41200 6 vssd1.extra22
port 712 nsew ground bidirectional
rlabel metal4 s 342804 -1864 343404 41200 6 vssd1.extra23
port 713 nsew ground bidirectional
rlabel metal4 s 306804 -1864 307404 41200 6 vssd1.extra24
port 714 nsew ground bidirectional
rlabel metal4 s 270804 -1864 271404 41200 6 vssd1.extra25
port 715 nsew ground bidirectional
rlabel metal4 s 234804 -1864 235404 41200 6 vssd1.extra26
port 716 nsew ground bidirectional
rlabel metal4 s 198804 -1864 199404 41200 6 vssd1.extra27
port 717 nsew ground bidirectional
rlabel metal4 s 162804 -1864 163404 41200 6 vssd1.extra28
port 718 nsew ground bidirectional
rlabel metal4 s 126804 -1864 127404 41200 6 vssd1.extra29
port 719 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 41200 6 vssd1.extra30
port 720 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1.extra31
port 721 nsew ground bidirectional
rlabel metal5 s -2936 667876 586860 668476 6 vssd1.extra32
port 722 nsew ground bidirectional
rlabel metal5 s -2936 631876 586860 632476 6 vssd1.extra33
port 723 nsew ground bidirectional
rlabel metal5 s -2936 595876 586860 596476 6 vssd1.extra34
port 724 nsew ground bidirectional
rlabel metal5 s -2936 559876 586860 560476 6 vssd1.extra35
port 725 nsew ground bidirectional
rlabel metal5 s -2936 523876 586860 524476 6 vssd1.extra36
port 726 nsew ground bidirectional
rlabel metal5 s -2936 487876 586860 488476 6 vssd1.extra37
port 727 nsew ground bidirectional
rlabel metal5 s -2936 451876 586860 452476 6 vssd1.extra38
port 728 nsew ground bidirectional
rlabel metal5 s -2936 415876 586860 416476 6 vssd1.extra39
port 729 nsew ground bidirectional
rlabel metal5 s -2936 379876 586860 380476 6 vssd1.extra40
port 730 nsew ground bidirectional
rlabel metal5 s -2936 343876 586860 344476 6 vssd1.extra41
port 731 nsew ground bidirectional
rlabel metal5 s -2936 307876 586860 308476 6 vssd1.extra42
port 732 nsew ground bidirectional
rlabel metal5 s -2936 271876 586860 272476 6 vssd1.extra43
port 733 nsew ground bidirectional
rlabel metal5 s -2936 235876 586860 236476 6 vssd1.extra44
port 734 nsew ground bidirectional
rlabel metal5 s -2936 199876 586860 200476 6 vssd1.extra45
port 735 nsew ground bidirectional
rlabel metal5 s -2936 163876 586860 164476 6 vssd1.extra46
port 736 nsew ground bidirectional
rlabel metal5 s -2936 127876 586860 128476 6 vssd1.extra47
port 737 nsew ground bidirectional
rlabel metal5 s -2936 91876 586860 92476 6 vssd1.extra48
port 738 nsew ground bidirectional
rlabel metal5 s -2936 55876 586860 56476 6 vssd1.extra49
port 739 nsew ground bidirectional
rlabel metal5 s -2936 19876 586860 20476 6 vssd1.extra50
port 740 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1.extra51
port 741 nsew ground bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 742 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2.extra1
port 743 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2.extra2
port 744 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2.extra3
port 745 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 746 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2.extra1
port 747 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2.extra2
port 748 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2.extra3
port 749 nsew ground bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 750 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1.extra1
port 751 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1.extra2
port 752 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1.extra3
port 753 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 754 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1.extra1
port 755 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1.extra2
port 756 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1.extra3
port 757 nsew ground bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 758 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2.extra1
port 759 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2.extra2
port 760 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2.extra3
port 761 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 762 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2.extra1
port 763 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2.extra2
port 764 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2.extra3
port 765 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
